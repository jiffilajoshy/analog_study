VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_vco_mix_dac
  CLASS BLOCK ;
  FOREIGN tt_um_vco_mix_dac ;
  ORIGIN -0.985 0.010 ;
  SIZE 152.090 BY 225.790 ;
  PIN inv_out_90
    ANTENNADIFFAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT 8.460 9.465 8.910 9.865 ;
    END
  END inv_out_90
  PIN inv_in_90
    ANTENNAGATEAREA 0.900000 ;
    ANTENNADIFFAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT 10.060 9.565 10.260 9.765 ;
    END
  END inv_in_90
  PIN inv_out_360
    ANTENNADIFFAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT 24.855 9.465 25.305 9.865 ;
    END
  END inv_out_360
  PIN inv_in_360
    ANTENNAGATEAREA 0.900000 ;
    ANTENNADIFFAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT 23.505 9.565 23.705 9.765 ;
    END
  END inv_in_360
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 63.345 119.165 63.945 123.165 ;
    END
  END clk
  PIN clk_out
    ANTENNAGATEAREA 1.140000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 87.145 119.165 87.745 123.165 ;
    END
  END clk_out
  PIN config[0]
    ANTENNAGATEAREA 263.660980 ;
    ANTENNADIFFAREA 130.662994 ;
    PORT
      LAYER met3 ;
        RECT 73.545 119.165 74.145 123.165 ;
    END
  END config[0]
  PIN config[10]
    ANTENNAGATEAREA 2.761500 ;
    PORT
      LAYER met3 ;
        RECT 83.745 119.165 84.345 123.165 ;
    END
  END config[10]
  PIN config[11]
    ANTENNAGATEAREA 2.439000 ;
    PORT
      LAYER met3 ;
        RECT 93.945 119.165 94.545 123.165 ;
    END
  END config[11]
  PIN config[1]
    ANTENNAGATEAREA 1.219500 ;
    PORT
      LAYER met3 ;
        RECT 97.345 119.165 97.945 123.165 ;
    END
  END config[1]
  PIN config[2]
    ANTENNAGATEAREA 260.576996 ;
    ANTENNADIFFAREA 130.662994 ;
    PORT
      LAYER met3 ;
        RECT 66.745 119.165 67.345 123.165 ;
    END
  END config[2]
  PIN config[3]
    ANTENNAGATEAREA 0.897000 ;
    PORT
      LAYER met3 ;
        RECT 80.345 119.165 80.945 123.165 ;
    END
  END config[3]
  PIN config[4]
    ANTENNAGATEAREA 0.967500 ;
    PORT
      LAYER met3 ;
        RECT 104.145 119.165 104.745 123.165 ;
    END
  END config[4]
  PIN config[5]
    ANTENNAGATEAREA 260.254486 ;
    ANTENNADIFFAREA 130.662994 ;
    PORT
      LAYER met3 ;
        RECT 70.145 119.165 70.745 123.165 ;
    END
  END config[5]
  PIN config[6]
    ANTENNAGATEAREA 0.322500 ;
    PORT
      LAYER met3 ;
        RECT 107.545 119.165 108.145 123.165 ;
    END
  END config[6]
  PIN config[7]
    ANTENNAGATEAREA 0.322500 ;
    PORT
      LAYER met3 ;
        RECT 76.945 119.165 77.545 123.165 ;
    END
  END config[7]
  PIN config[8]
    ANTENNAGATEAREA 0.322500 ;
    PORT
      LAYER met3 ;
        RECT 100.745 119.165 101.345 123.165 ;
    END
  END config[8]
  PIN config[9]
    ANTENNAGATEAREA 0.322500 ;
    PORT
      LAYER met3 ;
        RECT 90.545 119.165 91.145 123.165 ;
    END
  END config[9]
  PIN VGND
    ANTENNAGATEAREA 259.932007 ;
    ANTENNADIFFAREA 130.662994 ;
    PORT
      LAYER met4 ;
        RECT 60.345 96.625 112.505 98.625 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  PIN VPWR
    ANTENNAGATEAREA 164.229996 ;
    ANTENNADIFFAREA 188.643188 ;
    PORT
      LAYER met4 ;
        RECT 60.345 100.325 112.505 102.325 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT 16.115 202.035 17.825 203.295 ;
        RECT 19.265 202.035 20.975 203.295 ;
        RECT 23.040 202.040 24.750 203.300 ;
        RECT 27.430 202.045 29.140 203.305 ;
        RECT 31.685 202.040 33.395 203.300 ;
      LAYER nwell ;
        RECT 15.965 198.655 17.815 201.055 ;
        RECT 19.115 198.655 20.965 201.055 ;
        RECT 22.885 196.650 24.735 201.050 ;
        RECT 27.365 192.730 29.215 201.055 ;
        RECT 31.615 184.830 33.465 201.055 ;
      LAYER pwell ;
        RECT 60.690 117.500 61.500 117.640 ;
        RECT 60.500 117.330 61.500 117.500 ;
        RECT 60.690 116.270 61.500 117.330 ;
        RECT 60.690 116.120 61.500 116.260 ;
        RECT 60.500 115.950 61.500 116.120 ;
        RECT 60.690 113.510 61.500 115.950 ;
        RECT 60.690 113.360 61.370 113.500 ;
        RECT 60.500 113.190 61.370 113.360 ;
        RECT 60.690 109.985 61.370 113.190 ;
        RECT 60.690 109.075 61.590 109.985 ;
        RECT 60.690 107.540 61.370 109.075 ;
        RECT 60.690 105.770 61.600 107.540 ;
        RECT 60.535 105.370 60.645 105.530 ;
        RECT 60.775 104.320 61.560 104.750 ;
        RECT 60.690 104.160 61.500 104.300 ;
        RECT 60.500 103.990 61.500 104.160 ;
        RECT 60.690 98.790 61.500 103.990 ;
        RECT 60.535 98.470 60.645 98.630 ;
        RECT 60.690 97.715 61.600 97.860 ;
        RECT 60.500 97.545 61.600 97.715 ;
        RECT 60.690 95.670 61.600 97.545 ;
        RECT 60.690 95.420 61.500 95.560 ;
        RECT 60.500 95.250 61.500 95.420 ;
        RECT 60.690 91.890 61.500 95.250 ;
        RECT 60.775 91.440 61.560 91.870 ;
        RECT 60.690 89.445 61.600 91.320 ;
        RECT 60.500 89.275 61.600 89.445 ;
        RECT 60.690 89.130 61.600 89.275 ;
        RECT 60.690 88.980 61.500 89.120 ;
        RECT 60.500 88.810 61.500 88.980 ;
        RECT 60.690 83.610 61.500 88.810 ;
        RECT 60.690 83.460 61.500 83.600 ;
        RECT 60.500 83.290 61.500 83.460 ;
        RECT 60.690 82.230 61.500 83.290 ;
        RECT 60.690 82.075 61.370 82.220 ;
        RECT 60.500 81.905 61.370 82.075 ;
        RECT 60.690 80.375 61.370 81.905 ;
        RECT 60.690 79.010 61.600 80.375 ;
        RECT 60.775 78.560 61.560 78.990 ;
        RECT 60.690 78.400 61.500 78.540 ;
        RECT 60.500 78.230 61.500 78.400 ;
        RECT 60.690 73.030 61.500 78.230 ;
        RECT 60.690 72.880 61.500 73.020 ;
        RECT 60.500 72.710 61.500 72.880 ;
        RECT 60.690 67.510 61.500 72.710 ;
        RECT 60.530 67.245 60.640 67.365 ;
        RECT 60.690 65.980 61.500 67.040 ;
        RECT 60.500 65.810 61.500 65.980 ;
        RECT 60.690 65.670 61.500 65.810 ;
      LAYER nwell ;
        RECT 61.890 65.475 64.720 117.835 ;
      LAYER pwell ;
        RECT 65.110 117.500 65.920 117.640 ;
        RECT 66.130 117.500 66.940 117.640 ;
        RECT 65.110 117.330 66.940 117.500 ;
        RECT 65.110 116.270 65.920 117.330 ;
        RECT 66.130 116.270 66.940 117.330 ;
        RECT 65.110 116.120 65.920 116.260 ;
        RECT 66.130 116.120 66.940 116.260 ;
        RECT 65.110 115.950 66.940 116.120 ;
        RECT 65.110 113.510 65.920 115.950 ;
        RECT 66.130 114.430 66.940 115.950 ;
        RECT 65.970 114.165 66.080 114.285 ;
        RECT 66.130 113.810 66.910 113.960 ;
        RECT 65.940 113.640 66.910 113.810 ;
        RECT 65.240 113.360 65.920 113.500 ;
        RECT 65.240 113.190 66.110 113.360 ;
        RECT 65.240 109.985 65.920 113.190 ;
        RECT 66.130 112.590 66.910 113.640 ;
        RECT 66.130 112.440 66.810 112.580 ;
        RECT 65.940 112.270 66.810 112.440 ;
        RECT 65.020 109.075 65.920 109.985 ;
        RECT 65.240 107.540 65.920 109.075 ;
        RECT 65.010 105.770 65.920 107.540 ;
        RECT 66.130 109.065 66.810 112.270 ;
        RECT 66.130 108.155 67.030 109.065 ;
        RECT 66.130 106.620 66.810 108.155 ;
        RECT 65.110 105.540 65.920 105.680 ;
        RECT 65.110 105.370 66.110 105.540 ;
        RECT 65.110 103.850 65.920 105.370 ;
        RECT 66.130 104.850 67.040 106.620 ;
        RECT 66.215 104.320 67.000 104.750 ;
        RECT 65.975 103.990 66.085 104.150 ;
        RECT 65.010 102.455 65.920 103.825 ;
        RECT 66.160 103.235 66.840 103.380 ;
        RECT 65.940 103.065 66.840 103.235 ;
        RECT 65.240 101.865 65.920 102.455 ;
        RECT 65.240 101.695 66.110 101.865 ;
        RECT 65.240 101.550 65.920 101.695 ;
        RECT 66.160 101.575 66.840 103.065 ;
        RECT 65.010 95.880 65.920 101.390 ;
        RECT 66.130 100.175 67.040 101.575 ;
        RECT 65.970 99.905 66.080 100.025 ;
        RECT 66.130 96.500 66.810 99.470 ;
        RECT 66.130 96.155 67.040 96.500 ;
        RECT 65.940 95.985 67.040 96.155 ;
        RECT 65.010 95.710 66.110 95.880 ;
        RECT 65.010 95.570 65.920 95.710 ;
        RECT 66.130 95.570 67.040 95.985 ;
        RECT 65.110 95.420 65.920 95.560 ;
        RECT 65.970 95.420 66.080 95.425 ;
        RECT 65.110 95.250 66.110 95.420 ;
        RECT 65.110 94.190 65.920 95.250 ;
        RECT 65.010 92.795 65.920 94.165 ;
        RECT 66.130 93.705 67.040 95.100 ;
        RECT 65.240 92.205 65.920 92.795 ;
        RECT 66.160 93.690 67.040 93.705 ;
        RECT 66.160 92.660 66.840 93.690 ;
        RECT 65.940 92.490 66.840 92.660 ;
        RECT 66.160 92.365 66.840 92.490 ;
        RECT 65.240 92.035 66.110 92.205 ;
        RECT 65.240 91.890 65.920 92.035 ;
        RECT 65.050 91.440 65.835 91.870 ;
        RECT 65.110 91.280 65.920 91.420 ;
        RECT 65.110 91.110 66.110 91.280 ;
        RECT 65.110 89.590 65.920 91.110 ;
        RECT 65.240 89.440 65.920 89.580 ;
        RECT 65.240 89.270 66.110 89.440 ;
        RECT 65.240 86.065 65.920 89.270 ;
        RECT 66.130 88.985 67.040 92.270 ;
        RECT 65.940 88.815 67.040 88.985 ;
        RECT 66.130 88.670 67.040 88.815 ;
        RECT 65.020 85.155 65.920 86.065 ;
        RECT 66.130 85.765 67.040 88.660 ;
        RECT 65.940 85.620 67.040 85.765 ;
        RECT 65.940 85.595 66.110 85.620 ;
        RECT 66.130 85.300 66.940 85.440 ;
        RECT 65.240 83.620 65.920 85.155 ;
        RECT 65.940 85.130 66.940 85.300 ;
        RECT 66.130 84.070 66.940 85.130 ;
        RECT 66.130 83.915 66.810 84.060 ;
        RECT 65.940 83.745 66.810 83.915 ;
        RECT 65.010 81.850 65.920 83.620 ;
        RECT 66.130 81.980 66.810 83.745 ;
        RECT 65.240 81.620 65.920 81.760 ;
        RECT 65.240 81.450 66.110 81.620 ;
        RECT 65.240 78.245 65.920 81.450 ;
        RECT 66.130 80.390 67.040 81.980 ;
        RECT 66.130 80.240 66.940 80.380 ;
        RECT 65.940 80.070 66.940 80.240 ;
        RECT 66.130 79.010 66.940 80.070 ;
        RECT 66.215 78.560 67.000 78.990 ;
        RECT 66.130 78.400 66.940 78.540 ;
        RECT 65.020 77.335 65.920 78.245 ;
        RECT 65.940 78.230 66.940 78.400 ;
        RECT 65.240 75.800 65.920 77.335 ;
        RECT 65.010 74.030 65.920 75.800 ;
        RECT 65.110 73.800 65.920 73.940 ;
        RECT 65.110 73.630 66.110 73.800 ;
        RECT 65.110 68.430 65.920 73.630 ;
        RECT 66.130 73.030 66.940 78.230 ;
        RECT 66.130 72.880 66.940 73.020 ;
        RECT 65.940 72.710 66.940 72.880 ;
        RECT 65.110 68.280 65.920 68.420 ;
        RECT 65.110 68.110 66.110 68.280 ;
        RECT 65.110 67.050 65.920 68.110 ;
        RECT 66.130 67.510 66.940 72.710 ;
        RECT 65.970 67.245 66.080 67.365 ;
        RECT 65.110 65.980 65.920 67.040 ;
        RECT 66.130 65.980 66.940 67.040 ;
        RECT 65.110 65.810 66.940 65.980 ;
        RECT 65.110 65.670 65.920 65.810 ;
        RECT 66.130 65.670 66.940 65.810 ;
      LAYER nwell ;
        RECT 67.330 65.475 70.160 117.835 ;
      LAYER pwell ;
        RECT 70.550 117.500 71.360 117.640 ;
        RECT 71.570 117.500 72.380 117.640 ;
        RECT 70.550 117.330 72.380 117.500 ;
        RECT 70.550 116.270 71.360 117.330 ;
        RECT 71.570 116.270 72.380 117.330 ;
        RECT 70.550 116.120 71.360 116.260 ;
        RECT 71.410 116.120 71.520 116.125 ;
        RECT 70.550 115.950 71.550 116.120 ;
        RECT 70.550 114.890 71.360 115.950 ;
        RECT 71.800 115.655 72.480 115.800 ;
        RECT 71.380 115.485 72.480 115.655 ;
        RECT 70.650 114.735 71.330 114.880 ;
        RECT 70.650 114.565 71.550 114.735 ;
        RECT 70.650 113.075 71.330 114.565 ;
        RECT 70.450 111.675 71.360 113.075 ;
        RECT 71.570 112.600 72.480 115.485 ;
        RECT 71.570 112.440 72.250 112.580 ;
        RECT 71.380 112.270 72.250 112.440 ;
        RECT 70.580 111.510 71.360 111.660 ;
        RECT 70.580 111.340 71.550 111.510 ;
        RECT 70.580 110.290 71.360 111.340 ;
        RECT 70.550 110.140 71.360 110.280 ;
        RECT 70.550 109.970 71.550 110.140 ;
        RECT 70.550 106.610 71.360 109.970 ;
        RECT 71.570 109.065 72.250 112.270 ;
        RECT 71.570 108.155 72.470 109.065 ;
        RECT 71.570 106.620 72.250 108.155 ;
        RECT 70.450 106.465 71.360 106.590 ;
        RECT 70.450 106.295 71.550 106.465 ;
        RECT 70.450 103.390 71.360 106.295 ;
        RECT 71.570 104.850 72.480 106.620 ;
        RECT 71.655 104.320 72.440 104.750 ;
        RECT 71.570 104.160 72.380 104.300 ;
        RECT 71.380 103.990 72.380 104.160 ;
        RECT 70.450 100.025 71.360 103.360 ;
        RECT 71.570 102.470 72.380 103.990 ;
        RECT 71.410 102.205 71.520 102.325 ;
        RECT 71.570 101.860 72.480 102.000 ;
        RECT 71.380 101.690 72.480 101.860 ;
        RECT 70.450 99.855 71.550 100.025 ;
        RECT 70.450 99.710 71.360 99.855 ;
        RECT 70.550 99.560 71.360 99.700 ;
        RECT 70.550 99.390 71.550 99.560 ;
        RECT 70.550 98.330 71.360 99.390 ;
        RECT 70.450 98.180 71.360 98.320 ;
        RECT 70.450 98.010 71.550 98.180 ;
        RECT 70.450 95.110 71.360 98.010 ;
        RECT 71.570 96.180 72.480 101.690 ;
        RECT 70.650 94.960 71.330 95.085 ;
        RECT 70.650 94.790 71.550 94.960 ;
        RECT 70.650 93.760 71.330 94.790 ;
        RECT 70.450 92.380 71.360 93.760 ;
        RECT 71.410 92.085 71.520 92.205 ;
        RECT 70.490 91.440 71.275 91.870 ;
        RECT 70.550 91.280 71.360 91.420 ;
        RECT 70.550 91.110 71.550 91.280 ;
        RECT 70.550 90.050 71.360 91.110 ;
        RECT 70.680 89.900 71.360 90.040 ;
        RECT 70.680 89.730 71.550 89.900 ;
        RECT 70.680 86.525 71.360 89.730 ;
        RECT 71.570 87.140 72.250 95.935 ;
        RECT 71.380 86.970 72.250 87.140 ;
        RECT 71.570 86.830 72.250 86.970 ;
        RECT 70.460 85.615 71.360 86.525 ;
        RECT 70.680 84.080 71.360 85.615 ;
        RECT 71.570 85.425 72.480 86.820 ;
        RECT 71.600 85.410 72.480 85.425 ;
        RECT 71.600 84.380 72.280 85.410 ;
        RECT 71.380 84.210 72.280 84.380 ;
        RECT 71.600 84.085 72.280 84.210 ;
        RECT 70.450 82.310 71.360 84.080 ;
        RECT 71.410 83.805 71.520 83.925 ;
        RECT 70.450 80.370 71.360 82.140 ;
        RECT 71.570 80.705 72.480 83.600 ;
        RECT 71.380 80.535 72.480 80.705 ;
        RECT 71.570 80.390 72.480 80.535 ;
        RECT 70.680 78.835 71.360 80.370 ;
        RECT 71.570 80.240 72.480 80.370 ;
        RECT 71.380 80.070 72.480 80.240 ;
        RECT 71.570 79.020 72.480 80.070 ;
        RECT 70.460 77.925 71.360 78.835 ;
        RECT 71.655 78.560 72.440 78.990 ;
        RECT 71.570 78.400 72.380 78.540 ;
        RECT 71.380 78.230 72.380 78.400 ;
        RECT 70.680 74.720 71.360 77.925 ;
        RECT 70.680 74.550 71.550 74.720 ;
        RECT 70.680 74.410 71.360 74.550 ;
        RECT 70.650 74.260 71.330 74.385 ;
        RECT 70.650 74.090 71.550 74.260 ;
        RECT 70.650 73.060 71.330 74.090 ;
        RECT 70.450 73.045 71.330 73.060 ;
        RECT 70.450 71.650 71.360 73.045 ;
        RECT 71.570 73.030 72.380 78.230 ;
        RECT 71.570 72.880 72.380 73.020 ;
        RECT 71.380 72.710 72.380 72.880 ;
        RECT 70.550 71.500 71.360 71.640 ;
        RECT 70.550 71.330 71.550 71.500 ;
        RECT 70.550 67.970 71.360 71.330 ;
        RECT 71.405 67.650 71.515 67.810 ;
        RECT 71.570 67.510 72.380 72.710 ;
        RECT 71.410 67.245 71.520 67.365 ;
        RECT 70.550 65.980 71.360 67.040 ;
        RECT 71.570 65.980 72.380 67.040 ;
        RECT 70.550 65.810 72.380 65.980 ;
        RECT 70.550 65.670 71.360 65.810 ;
        RECT 71.570 65.670 72.380 65.810 ;
      LAYER nwell ;
        RECT 72.770 65.475 75.600 117.835 ;
      LAYER pwell ;
        RECT 75.990 117.500 76.800 117.640 ;
        RECT 77.010 117.500 77.820 117.640 ;
        RECT 75.990 117.330 77.820 117.500 ;
        RECT 75.990 116.270 76.800 117.330 ;
        RECT 77.010 116.270 77.820 117.330 ;
        RECT 75.990 116.120 76.800 116.260 ;
        RECT 77.010 116.120 77.820 116.260 ;
        RECT 75.990 115.950 77.820 116.120 ;
        RECT 75.990 114.890 76.800 115.950 ;
        RECT 77.010 114.890 77.820 115.950 ;
        RECT 75.890 114.735 76.570 114.880 ;
        RECT 77.040 114.735 77.720 114.880 ;
        RECT 75.890 114.565 77.720 114.735 ;
        RECT 75.890 111.680 76.800 114.565 ;
        RECT 77.040 113.075 77.720 114.565 ;
        RECT 77.010 111.675 77.920 113.075 ;
        RECT 76.090 111.520 76.770 111.645 ;
        RECT 77.010 111.520 77.820 111.660 ;
        RECT 76.090 111.350 77.820 111.520 ;
        RECT 76.090 110.320 76.770 111.350 ;
        RECT 75.890 108.940 76.800 110.320 ;
        RECT 75.990 108.760 76.800 108.900 ;
        RECT 75.990 108.590 76.990 108.760 ;
        RECT 75.990 103.390 76.800 108.590 ;
        RECT 77.010 106.150 77.820 111.350 ;
        RECT 77.010 106.000 77.820 106.140 ;
        RECT 76.820 105.830 77.820 106.000 ;
        RECT 77.010 104.770 77.820 105.830 ;
        RECT 77.095 104.320 77.880 104.750 ;
        RECT 77.010 104.160 77.820 104.300 ;
        RECT 76.820 103.990 77.820 104.160 ;
        RECT 75.990 103.240 76.800 103.380 ;
        RECT 75.990 103.070 76.990 103.240 ;
        RECT 75.990 97.870 76.800 103.070 ;
        RECT 77.010 98.790 77.820 103.990 ;
        RECT 77.010 98.640 77.820 98.780 ;
        RECT 76.820 98.470 77.820 98.640 ;
        RECT 75.990 97.720 76.800 97.860 ;
        RECT 75.990 97.550 76.990 97.720 ;
        RECT 75.990 92.350 76.800 97.550 ;
        RECT 77.010 93.270 77.820 98.470 ;
        RECT 76.855 92.950 76.965 93.110 ;
        RECT 76.850 92.200 76.960 92.205 ;
        RECT 77.010 92.200 77.920 92.340 ;
        RECT 76.820 92.030 77.920 92.200 ;
        RECT 75.930 91.440 76.715 91.870 ;
        RECT 75.890 90.025 76.800 91.420 ;
        RECT 75.890 90.010 76.770 90.025 ;
        RECT 76.090 88.980 76.770 90.010 ;
        RECT 76.090 88.810 76.990 88.980 ;
        RECT 76.090 88.685 76.770 88.810 ;
        RECT 75.990 88.520 76.800 88.660 ;
        RECT 75.990 88.350 76.990 88.520 ;
        RECT 75.990 83.150 76.800 88.350 ;
        RECT 77.010 86.500 77.920 92.030 ;
        RECT 77.010 86.220 77.820 86.360 ;
        RECT 76.820 86.050 77.820 86.220 ;
        RECT 75.990 83.000 76.800 83.140 ;
        RECT 75.990 82.830 76.990 83.000 ;
        RECT 75.990 81.310 76.800 82.830 ;
        RECT 77.010 82.690 77.820 86.050 ;
        RECT 76.855 82.370 76.965 82.530 ;
        RECT 77.040 81.620 77.720 81.745 ;
        RECT 76.820 81.450 77.720 81.620 ;
        RECT 75.890 79.915 76.800 81.285 ;
        RECT 77.040 80.420 77.720 81.450 ;
        RECT 77.040 80.405 77.920 80.420 ;
        RECT 76.120 79.325 76.800 79.915 ;
        RECT 76.120 79.155 76.990 79.325 ;
        RECT 76.120 79.010 76.800 79.155 ;
        RECT 77.010 79.010 77.920 80.405 ;
        RECT 75.990 78.860 76.800 79.000 ;
        RECT 75.990 78.690 76.990 78.860 ;
        RECT 75.990 73.490 76.800 78.690 ;
        RECT 77.095 78.560 77.880 78.990 ;
        RECT 77.010 78.400 77.690 78.540 ;
        RECT 76.820 78.230 77.690 78.400 ;
        RECT 77.010 75.025 77.690 78.230 ;
        RECT 77.010 74.115 77.910 75.025 ;
        RECT 75.990 73.340 76.800 73.480 ;
        RECT 75.990 73.170 76.990 73.340 ;
        RECT 75.990 67.970 76.800 73.170 ;
        RECT 77.010 72.580 77.690 74.115 ;
        RECT 77.010 70.810 77.920 72.580 ;
        RECT 77.010 70.580 77.820 70.720 ;
        RECT 76.820 70.410 77.820 70.580 ;
        RECT 76.845 67.650 76.955 67.810 ;
        RECT 77.010 67.050 77.820 70.410 ;
        RECT 75.990 65.980 76.800 67.040 ;
        RECT 77.010 65.980 77.820 67.040 ;
        RECT 75.990 65.810 77.820 65.980 ;
        RECT 75.990 65.670 76.800 65.810 ;
        RECT 77.010 65.670 77.820 65.810 ;
      LAYER nwell ;
        RECT 78.210 65.475 81.040 117.835 ;
      LAYER pwell ;
        RECT 81.430 117.500 82.240 117.640 ;
        RECT 82.450 117.500 83.260 117.640 ;
        RECT 81.430 117.330 83.260 117.500 ;
        RECT 81.430 116.270 82.240 117.330 ;
        RECT 82.450 116.270 83.260 117.330 ;
        RECT 81.460 116.110 82.240 116.260 ;
        RECT 82.450 116.120 83.260 116.260 ;
        RECT 82.260 116.110 83.260 116.120 ;
        RECT 81.460 115.950 83.260 116.110 ;
        RECT 81.460 115.940 82.430 115.950 ;
        RECT 81.460 114.890 82.240 115.940 ;
        RECT 81.460 114.730 82.240 114.880 ;
        RECT 81.460 114.560 82.430 114.730 ;
        RECT 81.460 113.510 82.240 114.560 ;
        RECT 82.450 114.430 83.260 115.950 ;
        RECT 82.290 114.165 82.400 114.285 ;
        RECT 82.450 113.820 83.130 113.960 ;
        RECT 82.260 113.650 83.130 113.820 ;
        RECT 81.560 113.360 82.240 113.500 ;
        RECT 81.560 113.190 82.430 113.360 ;
        RECT 81.560 109.985 82.240 113.190 ;
        RECT 81.340 109.075 82.240 109.985 ;
        RECT 81.560 107.540 82.240 109.075 ;
        RECT 81.330 105.770 82.240 107.540 ;
        RECT 82.450 110.445 83.130 113.650 ;
        RECT 82.450 109.535 83.350 110.445 ;
        RECT 82.450 108.000 83.130 109.535 ;
        RECT 82.450 106.230 83.360 108.000 ;
        RECT 82.450 106.000 83.260 106.140 ;
        RECT 82.260 105.830 83.260 106.000 ;
        RECT 82.285 105.370 82.395 105.530 ;
        RECT 82.450 104.770 83.260 105.830 ;
        RECT 81.330 103.350 82.240 104.730 ;
        RECT 82.535 104.320 83.320 104.750 ;
        RECT 82.295 103.990 82.405 104.150 ;
        RECT 81.530 102.320 82.210 103.350 ;
        RECT 81.530 102.150 82.430 102.320 ;
        RECT 81.530 102.025 82.210 102.150 ;
        RECT 81.330 101.860 82.240 102.000 ;
        RECT 81.330 101.690 82.430 101.860 ;
        RECT 81.330 96.180 82.240 101.690 ;
        RECT 82.450 100.475 83.360 103.380 ;
        RECT 82.260 100.305 83.360 100.475 ;
        RECT 82.450 100.180 83.360 100.305 ;
        RECT 82.450 100.020 83.260 100.160 ;
        RECT 82.260 99.850 83.260 100.020 ;
        RECT 82.450 98.790 83.260 99.850 ;
        RECT 82.450 98.640 83.360 98.690 ;
        RECT 82.260 98.470 83.360 98.640 ;
        RECT 81.330 94.625 82.240 96.020 ;
        RECT 81.330 94.610 82.210 94.625 ;
        RECT 81.530 93.580 82.210 94.610 ;
        RECT 82.450 94.200 83.360 98.470 ;
        RECT 82.295 93.870 82.405 94.030 ;
        RECT 81.530 93.410 82.430 93.580 ;
        RECT 81.530 93.285 82.210 93.410 ;
        RECT 81.430 93.120 82.240 93.260 ;
        RECT 82.450 93.120 83.360 93.260 ;
        RECT 81.430 92.950 83.360 93.120 ;
        RECT 81.430 91.890 82.240 92.950 ;
        RECT 81.370 91.440 82.155 91.870 ;
        RECT 81.330 89.570 82.240 91.340 ;
        RECT 81.560 88.035 82.240 89.570 ;
        RECT 81.340 87.125 82.240 88.035 ;
        RECT 82.450 87.420 83.360 92.950 ;
        RECT 82.450 87.140 83.260 87.280 ;
        RECT 81.560 83.920 82.240 87.125 ;
        RECT 82.260 86.970 83.260 87.140 ;
        RECT 81.560 83.750 82.430 83.920 ;
        RECT 81.560 83.610 82.240 83.750 ;
        RECT 82.450 83.610 83.260 86.970 ;
        RECT 81.430 83.460 82.240 83.600 ;
        RECT 82.450 83.460 83.260 83.600 ;
        RECT 81.430 83.290 83.260 83.460 ;
        RECT 81.430 81.770 82.240 83.290 ;
        RECT 82.450 82.230 83.260 83.290 ;
        RECT 82.290 81.505 82.400 81.625 ;
        RECT 81.530 81.160 82.210 81.285 ;
        RECT 81.530 80.990 82.430 81.160 ;
        RECT 81.530 79.960 82.210 80.990 ;
        RECT 81.330 79.945 82.210 79.960 ;
        RECT 81.330 78.550 82.240 79.945 ;
        RECT 82.450 79.325 83.360 82.220 ;
        RECT 82.260 79.180 83.360 79.325 ;
        RECT 82.260 79.155 82.430 79.180 ;
        RECT 82.535 78.560 83.320 78.990 ;
        RECT 81.330 78.395 82.240 78.540 ;
        RECT 82.290 78.395 82.400 78.405 ;
        RECT 81.330 78.225 82.430 78.395 ;
        RECT 81.330 76.350 82.240 78.225 ;
        RECT 82.450 77.940 83.130 78.080 ;
        RECT 82.260 77.770 83.130 77.940 ;
        RECT 81.430 76.100 82.240 76.240 ;
        RECT 81.430 75.930 82.430 76.100 ;
        RECT 81.430 70.730 82.240 75.930 ;
        RECT 82.450 74.565 83.130 77.770 ;
        RECT 82.450 73.655 83.350 74.565 ;
        RECT 82.450 72.120 83.130 73.655 ;
        RECT 81.430 70.580 82.240 70.720 ;
        RECT 81.430 70.410 82.430 70.580 ;
        RECT 81.430 67.050 82.240 70.410 ;
        RECT 82.450 70.350 83.360 72.120 ;
        RECT 82.450 70.120 83.260 70.260 ;
        RECT 82.260 69.950 83.260 70.120 ;
        RECT 82.450 67.510 83.260 69.950 ;
        RECT 82.290 67.245 82.400 67.365 ;
        RECT 81.430 65.980 82.240 67.040 ;
        RECT 82.450 65.980 83.260 67.040 ;
        RECT 81.430 65.810 83.260 65.980 ;
        RECT 81.430 65.670 82.240 65.810 ;
        RECT 82.450 65.670 83.260 65.810 ;
      LAYER nwell ;
        RECT 83.650 65.475 86.480 117.835 ;
      LAYER pwell ;
        RECT 86.870 117.500 87.680 117.640 ;
        RECT 87.890 117.500 88.700 117.640 ;
        RECT 86.870 117.330 88.700 117.500 ;
        RECT 86.870 116.270 87.680 117.330 ;
        RECT 87.890 116.270 88.700 117.330 ;
        RECT 86.870 116.120 87.680 116.260 ;
        RECT 86.870 116.110 87.870 116.120 ;
        RECT 87.890 116.110 88.670 116.260 ;
        RECT 86.870 115.950 88.670 116.110 ;
        RECT 86.870 110.750 87.680 115.950 ;
        RECT 87.700 115.940 88.670 115.950 ;
        RECT 87.890 114.890 88.670 115.940 ;
        RECT 87.890 114.740 88.570 114.880 ;
        RECT 87.700 114.570 88.570 114.740 ;
        RECT 87.890 111.365 88.570 114.570 ;
        RECT 86.870 110.600 87.680 110.740 ;
        RECT 86.870 110.430 87.870 110.600 ;
        RECT 87.890 110.455 88.790 111.365 ;
        RECT 86.870 107.070 87.680 110.430 ;
        RECT 87.890 108.920 88.570 110.455 ;
        RECT 87.890 107.150 88.800 108.920 ;
        RECT 87.730 106.920 87.840 106.925 ;
        RECT 87.890 106.920 88.700 107.060 ;
        RECT 87.700 106.750 88.700 106.920 ;
        RECT 86.970 106.455 87.650 106.600 ;
        RECT 86.970 106.285 87.870 106.455 ;
        RECT 86.970 104.795 87.650 106.285 ;
        RECT 87.890 105.230 88.700 106.750 ;
        RECT 87.730 104.965 87.840 105.085 ;
        RECT 86.770 103.395 87.680 104.795 ;
        RECT 87.975 104.320 88.760 104.750 ;
        RECT 87.890 104.155 88.800 104.300 ;
        RECT 87.700 103.985 88.800 104.155 ;
        RECT 86.770 103.235 87.680 103.380 ;
        RECT 86.770 103.065 87.870 103.235 ;
        RECT 86.770 100.170 87.680 103.065 ;
        RECT 86.770 100.020 87.680 100.160 ;
        RECT 86.770 99.850 87.870 100.020 ;
        RECT 86.770 96.950 87.680 99.850 ;
        RECT 87.890 99.750 88.800 103.985 ;
        RECT 87.730 99.445 87.840 99.565 ;
        RECT 87.890 99.100 88.800 99.240 ;
        RECT 87.700 98.930 88.800 99.100 ;
        RECT 86.970 96.795 87.650 96.940 ;
        RECT 86.970 96.625 87.870 96.795 ;
        RECT 86.970 95.135 87.650 96.625 ;
        RECT 87.890 96.030 88.800 98.930 ;
        RECT 87.920 95.875 88.600 96.020 ;
        RECT 87.700 95.705 88.600 95.875 ;
        RECT 86.770 93.735 87.680 95.135 ;
        RECT 87.920 94.215 88.600 95.705 ;
        RECT 86.870 93.580 87.680 93.720 ;
        RECT 86.870 93.410 87.870 93.580 ;
        RECT 86.870 91.890 87.680 93.410 ;
        RECT 87.890 92.815 88.800 94.215 ;
        RECT 87.890 92.660 88.700 92.800 ;
        RECT 87.700 92.490 88.700 92.660 ;
        RECT 86.810 91.440 87.595 91.870 ;
        RECT 87.890 91.430 88.700 92.490 ;
        RECT 87.000 91.280 87.680 91.420 ;
        RECT 87.000 91.275 87.870 91.280 ;
        RECT 87.920 91.275 88.600 91.420 ;
        RECT 87.000 91.110 88.600 91.275 ;
        RECT 87.000 82.315 87.680 91.110 ;
        RECT 87.700 91.105 88.600 91.110 ;
        RECT 87.920 89.615 88.600 91.105 ;
        RECT 87.890 88.215 88.800 89.615 ;
        RECT 87.890 88.060 88.700 88.200 ;
        RECT 87.700 87.890 88.700 88.060 ;
        RECT 87.890 82.690 88.700 87.890 ;
        RECT 87.735 82.370 87.845 82.530 ;
        RECT 86.770 80.630 87.680 82.220 ;
        RECT 87.920 81.620 88.600 81.745 ;
        RECT 87.700 81.450 88.600 81.620 ;
        RECT 87.000 78.865 87.680 80.630 ;
        RECT 87.920 80.420 88.600 81.450 ;
        RECT 87.920 80.405 88.800 80.420 ;
        RECT 87.890 79.010 88.800 80.405 ;
        RECT 87.000 78.695 87.870 78.865 ;
        RECT 87.000 78.550 87.680 78.695 ;
        RECT 87.975 78.560 88.760 78.990 ;
        RECT 86.970 78.400 87.650 78.525 ;
        RECT 86.970 78.230 87.870 78.400 ;
        RECT 86.970 77.200 87.650 78.230 ;
        RECT 87.890 77.480 88.800 78.530 ;
        RECT 87.700 77.310 88.800 77.480 ;
        RECT 86.770 77.185 87.650 77.200 ;
        RECT 86.770 75.790 87.680 77.185 ;
        RECT 87.890 77.180 88.800 77.310 ;
        RECT 87.890 77.020 88.570 77.160 ;
        RECT 87.700 76.850 88.570 77.020 ;
        RECT 86.770 74.395 87.680 75.765 ;
        RECT 87.000 73.805 87.680 74.395 ;
        RECT 87.000 73.635 87.870 73.805 ;
        RECT 87.890 73.645 88.570 76.850 ;
        RECT 87.000 73.490 87.680 73.635 ;
        RECT 86.770 73.340 87.680 73.470 ;
        RECT 86.770 73.170 87.870 73.340 ;
        RECT 86.770 72.120 87.680 73.170 ;
        RECT 87.890 72.735 88.790 73.645 ;
        RECT 86.870 71.960 87.680 72.100 ;
        RECT 86.870 71.790 87.870 71.960 ;
        RECT 86.870 68.430 87.680 71.790 ;
        RECT 87.890 71.200 88.570 72.735 ;
        RECT 87.890 69.430 88.800 71.200 ;
        RECT 87.890 69.200 88.700 69.340 ;
        RECT 87.700 69.030 88.700 69.200 ;
        RECT 86.870 68.280 87.680 68.420 ;
        RECT 86.870 68.110 87.870 68.280 ;
        RECT 86.870 67.050 87.680 68.110 ;
        RECT 87.890 67.510 88.700 69.030 ;
        RECT 87.730 67.245 87.840 67.365 ;
        RECT 86.870 65.980 87.680 67.040 ;
        RECT 87.890 65.980 88.700 67.040 ;
        RECT 86.870 65.810 88.700 65.980 ;
        RECT 86.870 65.670 87.680 65.810 ;
        RECT 87.890 65.670 88.700 65.810 ;
      LAYER nwell ;
        RECT 89.090 65.475 91.920 117.835 ;
      LAYER pwell ;
        RECT 92.310 117.500 93.120 117.640 ;
        RECT 93.330 117.500 94.140 117.640 ;
        RECT 92.310 117.330 94.140 117.500 ;
        RECT 92.310 116.270 93.120 117.330 ;
        RECT 93.330 116.270 94.140 117.330 ;
        RECT 92.340 116.110 93.120 116.260 ;
        RECT 93.330 116.120 94.140 116.260 ;
        RECT 93.140 116.110 94.140 116.120 ;
        RECT 92.340 115.950 94.140 116.110 ;
        RECT 92.340 115.940 93.310 115.950 ;
        RECT 92.340 114.890 93.120 115.940 ;
        RECT 92.440 114.740 93.120 114.880 ;
        RECT 92.440 114.570 93.310 114.740 ;
        RECT 92.440 111.365 93.120 114.570 ;
        RECT 92.220 110.455 93.120 111.365 ;
        RECT 93.330 110.750 94.140 115.950 ;
        RECT 93.330 110.600 94.140 110.740 ;
        RECT 92.440 108.920 93.120 110.455 ;
        RECT 93.140 110.430 94.140 110.600 ;
        RECT 92.210 107.150 93.120 108.920 ;
        RECT 92.310 106.920 93.120 107.060 ;
        RECT 92.310 106.750 93.310 106.920 ;
        RECT 92.310 105.230 93.120 106.750 ;
        RECT 93.330 105.230 94.140 110.430 ;
        RECT 93.170 104.965 93.280 105.085 ;
        RECT 92.440 102.000 93.120 104.760 ;
        RECT 93.415 104.320 94.200 104.750 ;
        RECT 93.175 103.990 93.285 104.150 ;
        RECT 93.360 103.240 94.040 103.365 ;
        RECT 93.140 103.070 94.040 103.240 ;
        RECT 93.360 102.040 94.040 103.070 ;
        RECT 92.210 100.930 93.120 102.000 ;
        RECT 92.210 100.760 93.310 100.930 ;
        RECT 92.210 100.630 93.120 100.760 ;
        RECT 93.330 100.660 94.240 102.040 ;
        RECT 92.310 100.480 93.120 100.620 ;
        RECT 93.330 100.480 94.240 100.620 ;
        RECT 92.310 100.310 94.240 100.480 ;
        RECT 92.310 98.790 93.120 100.310 ;
        RECT 93.170 98.525 93.280 98.645 ;
        RECT 92.410 98.175 93.090 98.320 ;
        RECT 92.410 98.005 93.310 98.175 ;
        RECT 92.410 96.515 93.090 98.005 ;
        RECT 93.330 97.410 94.240 100.310 ;
        RECT 92.210 95.115 93.120 96.515 ;
        RECT 92.410 94.955 93.090 95.100 ;
        RECT 92.410 94.785 93.310 94.955 ;
        RECT 92.410 93.295 93.090 94.785 ;
        RECT 92.210 91.895 93.120 93.295 ;
        RECT 92.250 91.440 93.035 91.870 ;
        RECT 92.210 85.760 93.120 91.290 ;
        RECT 93.330 88.520 94.010 97.315 ;
        RECT 93.140 88.350 94.010 88.520 ;
        RECT 93.330 88.210 94.010 88.350 ;
        RECT 93.330 86.350 94.240 88.120 ;
        RECT 92.210 85.590 93.310 85.760 ;
        RECT 92.210 85.450 93.120 85.590 ;
        RECT 92.410 85.300 93.090 85.425 ;
        RECT 92.410 85.130 93.310 85.300 ;
        RECT 92.410 84.100 93.090 85.130 ;
        RECT 92.210 84.085 93.090 84.100 ;
        RECT 93.330 84.815 94.010 86.350 ;
        RECT 92.210 82.690 93.120 84.085 ;
        RECT 93.330 83.905 94.230 84.815 ;
        RECT 92.410 82.540 93.090 82.665 ;
        RECT 92.410 82.370 93.310 82.540 ;
        RECT 92.410 81.340 93.090 82.370 ;
        RECT 92.210 81.325 93.090 81.340 ;
        RECT 92.210 79.930 93.120 81.325 ;
        RECT 93.330 80.700 94.010 83.905 ;
        RECT 93.140 80.530 94.010 80.700 ;
        RECT 93.330 80.390 94.010 80.530 ;
        RECT 93.330 80.240 94.140 80.380 ;
        RECT 93.140 80.070 94.140 80.240 ;
        RECT 93.170 79.665 93.280 79.785 ;
        RECT 92.410 79.320 93.090 79.445 ;
        RECT 92.410 79.150 93.310 79.320 ;
        RECT 92.410 78.120 93.090 79.150 ;
        RECT 93.330 79.010 94.140 80.070 ;
        RECT 93.415 78.560 94.200 78.990 ;
        RECT 93.170 78.285 93.280 78.405 ;
        RECT 92.210 78.105 93.090 78.120 ;
        RECT 92.210 76.710 93.120 78.105 ;
        RECT 93.330 77.940 94.010 78.080 ;
        RECT 93.140 77.770 94.010 77.940 ;
        RECT 92.310 76.560 93.120 76.700 ;
        RECT 92.310 76.390 93.310 76.560 ;
        RECT 92.310 71.190 93.120 76.390 ;
        RECT 93.330 74.565 94.010 77.770 ;
        RECT 93.330 73.655 94.230 74.565 ;
        RECT 93.330 72.120 94.010 73.655 ;
        RECT 92.310 71.040 93.120 71.180 ;
        RECT 92.310 70.870 93.310 71.040 ;
        RECT 92.310 67.510 93.120 70.870 ;
        RECT 93.330 70.350 94.240 72.120 ;
        RECT 93.330 70.120 94.140 70.260 ;
        RECT 93.140 69.950 94.140 70.120 ;
        RECT 93.330 67.510 94.140 69.950 ;
        RECT 93.170 67.245 93.280 67.365 ;
        RECT 92.310 65.980 93.120 67.040 ;
        RECT 93.330 65.980 94.140 67.040 ;
        RECT 92.310 65.810 94.140 65.980 ;
        RECT 92.310 65.670 93.120 65.810 ;
        RECT 93.330 65.670 94.140 65.810 ;
      LAYER nwell ;
        RECT 94.530 65.475 97.360 117.835 ;
      LAYER pwell ;
        RECT 97.750 117.500 98.560 117.640 ;
        RECT 98.770 117.500 99.580 117.640 ;
        RECT 97.750 117.330 99.580 117.500 ;
        RECT 97.750 116.270 98.560 117.330 ;
        RECT 98.770 116.270 99.580 117.330 ;
        RECT 97.750 116.120 98.560 116.260 ;
        RECT 98.770 116.120 99.580 116.260 ;
        RECT 97.750 115.950 99.580 116.120 ;
        RECT 97.750 114.890 98.560 115.950 ;
        RECT 97.850 114.735 98.530 114.880 ;
        RECT 97.850 114.565 98.750 114.735 ;
        RECT 97.850 113.075 98.530 114.565 ;
        RECT 98.770 114.430 99.580 115.950 ;
        RECT 98.770 114.280 99.450 114.420 ;
        RECT 98.580 114.110 99.450 114.280 ;
        RECT 97.650 111.675 98.560 113.075 ;
        RECT 97.780 110.610 98.560 111.660 ;
        RECT 98.770 110.905 99.450 114.110 ;
        RECT 97.780 110.440 98.750 110.610 ;
        RECT 97.780 110.290 98.560 110.440 ;
        RECT 97.750 110.140 98.560 110.280 ;
        RECT 97.750 109.970 98.750 110.140 ;
        RECT 98.770 109.995 99.670 110.905 ;
        RECT 97.750 104.770 98.560 109.970 ;
        RECT 98.770 108.460 99.450 109.995 ;
        RECT 98.770 106.690 99.680 108.460 ;
        RECT 98.770 106.460 99.580 106.600 ;
        RECT 98.580 106.290 99.580 106.460 ;
        RECT 98.770 104.770 99.580 106.290 ;
        RECT 98.605 104.450 98.715 104.610 ;
        RECT 98.855 104.320 99.640 104.750 ;
        RECT 98.610 104.045 98.720 104.165 ;
        RECT 97.650 103.705 98.560 103.830 ;
        RECT 97.650 103.695 98.750 103.705 ;
        RECT 98.800 103.695 99.480 103.840 ;
        RECT 97.650 103.535 99.480 103.695 ;
        RECT 97.650 100.630 98.560 103.535 ;
        RECT 98.580 103.525 99.480 103.535 ;
        RECT 98.800 102.035 99.480 103.525 ;
        RECT 98.770 100.635 99.680 102.035 ;
        RECT 97.650 100.480 98.560 100.620 ;
        RECT 97.650 100.310 98.750 100.480 ;
        RECT 97.650 94.800 98.560 100.310 ;
        RECT 98.770 98.645 99.680 100.540 ;
        RECT 98.580 98.475 99.680 98.645 ;
        RECT 98.770 98.330 99.680 98.475 ;
        RECT 98.770 98.180 99.580 98.320 ;
        RECT 98.580 98.010 99.580 98.180 ;
        RECT 98.770 96.490 99.580 98.010 ;
        RECT 98.770 95.085 99.680 96.480 ;
        RECT 98.800 95.070 99.680 95.085 ;
        RECT 97.880 94.500 98.560 94.640 ;
        RECT 97.880 94.330 98.750 94.500 ;
        RECT 97.880 91.900 98.560 94.330 ;
        RECT 98.800 94.040 99.480 95.070 ;
        RECT 98.580 93.870 99.480 94.040 ;
        RECT 98.800 93.745 99.480 93.870 ;
        RECT 98.770 93.580 99.580 93.720 ;
        RECT 98.580 93.410 99.580 93.580 ;
        RECT 97.690 91.440 98.475 91.870 ;
        RECT 97.650 89.445 98.560 91.340 ;
        RECT 97.650 89.275 98.750 89.445 ;
        RECT 97.650 89.130 98.560 89.275 ;
        RECT 97.750 88.980 98.560 89.120 ;
        RECT 97.750 88.810 98.750 88.980 ;
        RECT 97.750 86.370 98.560 88.810 ;
        RECT 98.770 88.210 99.580 93.410 ;
        RECT 98.770 88.060 99.580 88.200 ;
        RECT 98.580 87.890 99.580 88.060 ;
        RECT 98.610 86.105 98.720 86.225 ;
        RECT 98.580 85.730 98.750 85.755 ;
        RECT 97.650 85.585 98.750 85.730 ;
        RECT 97.650 82.690 98.560 85.585 ;
        RECT 98.770 82.690 99.580 87.890 ;
        RECT 97.650 81.620 98.560 82.670 ;
        RECT 98.610 82.425 98.720 82.545 ;
        RECT 97.650 81.450 98.750 81.620 ;
        RECT 97.650 81.320 98.560 81.450 ;
        RECT 97.750 81.160 98.560 81.300 ;
        RECT 97.750 80.990 98.750 81.160 ;
        RECT 97.750 79.470 98.560 80.990 ;
        RECT 98.770 80.825 99.680 82.220 ;
        RECT 98.800 80.810 99.680 80.825 ;
        RECT 98.800 79.780 99.480 80.810 ;
        RECT 98.580 79.610 99.480 79.780 ;
        RECT 98.800 79.485 99.480 79.610 ;
        RECT 97.650 77.485 98.560 79.360 ;
        RECT 98.610 79.205 98.720 79.325 ;
        RECT 98.855 78.560 99.640 78.990 ;
        RECT 97.650 77.315 98.750 77.485 ;
        RECT 97.650 77.170 98.560 77.315 ;
        RECT 97.880 77.015 98.560 77.160 ;
        RECT 98.770 77.155 99.680 78.525 ;
        RECT 97.880 76.845 98.750 77.015 ;
        RECT 97.880 76.255 98.560 76.845 ;
        RECT 98.770 76.565 99.450 77.155 ;
        RECT 98.580 76.395 99.450 76.565 ;
        RECT 97.650 74.885 98.560 76.255 ;
        RECT 98.770 76.250 99.450 76.395 ;
        RECT 98.770 76.100 99.580 76.240 ;
        RECT 98.580 75.930 99.580 76.100 ;
        RECT 97.750 74.720 98.560 74.860 ;
        RECT 97.750 74.550 98.750 74.720 ;
        RECT 97.750 69.350 98.560 74.550 ;
        RECT 98.770 70.730 99.580 75.930 ;
        RECT 98.770 70.580 99.580 70.720 ;
        RECT 98.580 70.410 99.580 70.580 ;
        RECT 97.750 69.200 98.560 69.340 ;
        RECT 97.750 69.030 98.750 69.200 ;
        RECT 97.750 67.510 98.560 69.030 ;
        RECT 98.610 67.245 98.720 67.365 ;
        RECT 98.770 67.050 99.580 70.410 ;
        RECT 97.750 65.980 98.560 67.040 ;
        RECT 98.770 65.980 99.580 67.040 ;
        RECT 97.750 65.810 99.580 65.980 ;
        RECT 97.750 65.670 98.560 65.810 ;
        RECT 98.770 65.670 99.580 65.810 ;
      LAYER nwell ;
        RECT 99.970 65.475 102.800 117.835 ;
      LAYER pwell ;
        RECT 103.190 117.500 104.000 117.640 ;
        RECT 104.210 117.500 105.020 117.640 ;
        RECT 103.190 117.330 105.020 117.500 ;
        RECT 103.190 116.270 104.000 117.330 ;
        RECT 104.210 116.270 105.020 117.330 ;
        RECT 103.220 116.110 104.000 116.260 ;
        RECT 103.220 115.940 104.190 116.110 ;
        RECT 103.220 114.890 104.000 115.940 ;
        RECT 104.210 115.190 104.990 115.340 ;
        RECT 104.020 115.020 104.990 115.190 ;
        RECT 103.220 114.730 104.000 114.880 ;
        RECT 103.220 114.560 104.190 114.730 ;
        RECT 103.220 113.510 104.000 114.560 ;
        RECT 104.210 113.970 104.990 115.020 ;
        RECT 104.210 113.820 104.890 113.960 ;
        RECT 104.020 113.650 104.890 113.820 ;
        RECT 103.320 113.360 104.000 113.500 ;
        RECT 103.320 113.190 104.190 113.360 ;
        RECT 103.320 109.985 104.000 113.190 ;
        RECT 103.100 109.075 104.000 109.985 ;
        RECT 103.320 107.540 104.000 109.075 ;
        RECT 103.090 105.770 104.000 107.540 ;
        RECT 104.210 110.445 104.890 113.650 ;
        RECT 104.210 109.535 105.110 110.445 ;
        RECT 104.210 108.000 104.890 109.535 ;
        RECT 104.210 106.230 105.120 108.000 ;
        RECT 104.210 106.000 105.020 106.140 ;
        RECT 104.020 105.830 105.020 106.000 ;
        RECT 104.050 105.425 104.160 105.545 ;
        RECT 103.320 105.075 104.000 105.220 ;
        RECT 103.320 104.905 104.190 105.075 ;
        RECT 103.320 104.315 104.000 104.905 ;
        RECT 104.210 104.770 105.020 105.830 ;
        RECT 104.295 104.320 105.080 104.750 ;
        RECT 103.090 102.945 104.000 104.315 ;
        RECT 104.210 104.160 105.020 104.300 ;
        RECT 104.020 103.990 105.020 104.160 ;
        RECT 104.210 102.930 105.020 103.990 ;
        RECT 104.210 102.780 105.120 102.920 ;
        RECT 104.020 102.610 105.120 102.780 ;
        RECT 103.090 101.855 104.000 102.000 ;
        RECT 103.090 101.685 104.190 101.855 ;
        RECT 103.090 99.790 104.000 101.685 ;
        RECT 103.190 99.560 104.000 99.700 ;
        RECT 103.190 99.390 104.190 99.560 ;
        RECT 103.190 97.870 104.000 99.390 ;
        RECT 103.090 97.720 104.000 97.860 ;
        RECT 103.090 97.550 104.190 97.720 ;
        RECT 103.090 92.020 104.000 97.550 ;
        RECT 104.210 97.080 105.120 102.610 ;
        RECT 104.050 96.685 104.160 96.805 ;
        RECT 104.210 94.630 105.120 96.400 ;
        RECT 104.210 93.095 104.890 94.630 ;
        RECT 104.210 92.185 105.110 93.095 ;
        RECT 103.130 91.440 103.915 91.870 ;
        RECT 103.090 85.760 104.000 91.290 ;
        RECT 104.210 88.980 104.890 92.185 ;
        RECT 104.020 88.810 104.890 88.980 ;
        RECT 104.210 88.670 104.890 88.810 ;
        RECT 104.210 88.520 105.020 88.660 ;
        RECT 104.020 88.350 105.020 88.520 ;
        RECT 104.210 86.830 105.020 88.350 ;
        RECT 104.210 86.680 104.890 86.820 ;
        RECT 104.020 86.510 104.890 86.680 ;
        RECT 103.090 85.590 104.190 85.760 ;
        RECT 103.090 85.450 104.000 85.590 ;
        RECT 104.020 85.270 104.190 85.300 ;
        RECT 103.180 85.130 104.190 85.270 ;
        RECT 103.180 84.290 104.000 85.130 ;
        RECT 103.090 82.700 104.000 84.290 ;
        RECT 104.210 83.305 104.890 86.510 ;
        RECT 104.050 82.425 104.160 82.545 ;
        RECT 104.210 82.395 105.110 83.305 ;
        RECT 103.320 82.080 104.000 82.220 ;
        RECT 103.320 81.910 104.190 82.080 ;
        RECT 103.320 78.705 104.000 81.910 ;
        RECT 104.210 80.860 104.890 82.395 ;
        RECT 104.210 79.090 105.120 80.860 ;
        RECT 103.100 77.795 104.000 78.705 ;
        RECT 104.295 78.560 105.080 78.990 ;
        RECT 104.210 78.395 105.120 78.540 ;
        RECT 104.020 78.225 105.120 78.395 ;
        RECT 103.320 76.260 104.000 77.795 ;
        RECT 104.210 76.350 105.120 78.225 ;
        RECT 103.090 74.490 104.000 76.260 ;
        RECT 104.210 76.100 105.020 76.240 ;
        RECT 104.020 75.930 105.020 76.100 ;
        RECT 103.090 74.255 104.000 74.400 ;
        RECT 103.090 74.085 104.190 74.255 ;
        RECT 103.090 72.210 104.000 74.085 ;
        RECT 103.190 71.960 104.000 72.100 ;
        RECT 103.190 71.790 104.190 71.960 ;
        RECT 103.190 68.430 104.000 71.790 ;
        RECT 104.210 70.730 105.020 75.930 ;
        RECT 104.210 70.580 105.020 70.720 ;
        RECT 104.020 70.410 105.020 70.580 ;
        RECT 103.190 68.280 104.000 68.420 ;
        RECT 103.190 68.110 104.190 68.280 ;
        RECT 103.190 67.050 104.000 68.110 ;
        RECT 104.210 67.050 105.020 70.410 ;
        RECT 103.190 65.980 104.000 67.040 ;
        RECT 104.210 65.980 105.020 67.040 ;
        RECT 103.190 65.810 105.020 65.980 ;
        RECT 103.190 65.670 104.000 65.810 ;
        RECT 104.210 65.670 105.020 65.810 ;
      LAYER nwell ;
        RECT 105.410 65.475 108.240 117.835 ;
      LAYER pwell ;
        RECT 108.630 117.500 109.440 117.640 ;
        RECT 109.650 117.500 110.460 117.640 ;
        RECT 108.630 117.330 110.460 117.500 ;
        RECT 108.630 116.270 109.440 117.330 ;
        RECT 109.650 116.270 110.460 117.330 ;
        RECT 108.630 116.120 109.440 116.260 ;
        RECT 109.650 116.120 110.460 116.260 ;
        RECT 108.630 115.950 110.460 116.120 ;
        RECT 108.630 113.510 109.440 115.950 ;
        RECT 108.760 113.360 109.440 113.500 ;
        RECT 108.760 113.190 109.630 113.360 ;
        RECT 108.760 109.985 109.440 113.190 ;
        RECT 109.650 110.750 110.460 115.950 ;
        RECT 109.650 110.600 110.460 110.740 ;
        RECT 109.460 110.430 110.460 110.600 ;
        RECT 108.540 109.075 109.440 109.985 ;
        RECT 108.760 107.540 109.440 109.075 ;
        RECT 108.530 105.770 109.440 107.540 ;
        RECT 108.630 105.540 109.440 105.680 ;
        RECT 108.630 105.370 109.630 105.540 ;
        RECT 108.630 104.310 109.440 105.370 ;
        RECT 109.650 105.230 110.460 110.430 ;
        RECT 109.490 104.965 109.600 105.085 ;
        RECT 109.735 104.320 110.520 104.750 ;
        RECT 108.530 104.160 109.440 104.300 ;
        RECT 109.650 104.160 110.460 104.300 ;
        RECT 108.530 103.990 110.460 104.160 ;
        RECT 108.530 98.480 109.440 103.990 ;
        RECT 109.650 98.790 110.460 103.990 ;
        RECT 109.650 98.640 110.460 98.780 ;
        RECT 109.460 98.470 110.460 98.640 ;
        RECT 108.530 98.180 109.440 98.320 ;
        RECT 108.530 98.010 109.630 98.180 ;
        RECT 108.530 92.480 109.440 98.010 ;
        RECT 109.650 93.270 110.460 98.470 ;
        RECT 109.650 93.120 110.460 93.260 ;
        RECT 109.460 92.950 110.460 93.120 ;
        RECT 109.490 92.085 109.600 92.205 ;
        RECT 109.650 91.890 110.460 92.950 ;
        RECT 108.570 91.440 109.355 91.870 ;
        RECT 109.735 91.440 110.520 91.870 ;
        RECT 109.650 91.280 110.460 91.420 ;
        RECT 109.460 91.110 110.460 91.280 ;
        RECT 108.530 88.900 109.440 90.490 ;
        RECT 108.620 88.060 109.440 88.900 ;
        RECT 108.620 87.920 109.630 88.060 ;
        RECT 109.460 87.890 109.630 87.920 ;
        RECT 109.485 87.430 109.595 87.590 ;
        RECT 108.530 85.425 109.440 86.820 ;
        RECT 109.650 85.910 110.460 91.110 ;
        RECT 109.650 85.760 110.460 85.900 ;
        RECT 109.460 85.590 110.460 85.760 ;
        RECT 108.530 85.410 109.410 85.425 ;
        RECT 108.730 84.380 109.410 85.410 ;
        RECT 108.730 84.210 109.630 84.380 ;
        RECT 108.730 84.085 109.410 84.210 ;
        RECT 108.530 82.675 109.440 84.045 ;
        RECT 108.760 82.085 109.440 82.675 ;
        RECT 108.760 81.915 109.630 82.085 ;
        RECT 108.760 81.770 109.440 81.915 ;
        RECT 108.630 81.620 109.440 81.760 ;
        RECT 108.630 81.450 109.630 81.620 ;
        RECT 108.630 76.250 109.440 81.450 ;
        RECT 109.650 80.390 110.460 85.590 ;
        RECT 109.650 80.240 110.460 80.380 ;
        RECT 109.460 80.070 110.460 80.240 ;
        RECT 109.650 79.010 110.460 80.070 ;
        RECT 109.735 78.560 110.520 78.990 ;
        RECT 109.650 78.400 110.460 78.540 ;
        RECT 109.460 78.230 110.460 78.400 ;
        RECT 108.630 76.100 109.440 76.240 ;
        RECT 108.630 75.930 109.630 76.100 ;
        RECT 108.630 70.730 109.440 75.930 ;
        RECT 109.650 73.030 110.460 78.230 ;
        RECT 109.650 72.880 110.460 73.020 ;
        RECT 109.460 72.710 110.460 72.880 ;
        RECT 108.630 70.580 109.440 70.720 ;
        RECT 108.630 70.410 109.630 70.580 ;
        RECT 108.630 67.050 109.440 70.410 ;
        RECT 109.650 67.510 110.460 72.710 ;
        RECT 109.490 67.245 109.600 67.365 ;
        RECT 108.630 65.980 109.440 67.040 ;
        RECT 109.650 65.980 110.460 67.040 ;
        RECT 108.630 65.810 110.460 65.980 ;
        RECT 108.630 65.670 109.440 65.810 ;
        RECT 109.650 65.670 110.460 65.810 ;
      LAYER nwell ;
        RECT 110.850 65.475 112.455 117.835 ;
        RECT 12.225 19.470 14.075 21.870 ;
        RECT 15.845 19.475 17.695 21.875 ;
      LAYER pwell ;
        RECT 12.375 17.230 14.085 18.490 ;
        RECT 16.000 17.225 17.710 18.485 ;
        RECT 13.740 14.690 15.450 15.950 ;
        RECT 17.260 13.675 18.970 13.680 ;
        RECT 12.755 13.670 14.465 13.675 ;
        RECT 17.260 13.670 21.225 13.675 ;
        RECT 12.755 12.420 21.225 13.670 ;
        RECT 12.755 12.415 16.720 12.420 ;
        RECT 19.515 12.415 21.225 12.420 ;
        RECT 15.010 12.410 16.720 12.415 ;
        RECT 8.530 9.935 10.240 11.195 ;
        RECT 23.525 9.935 25.235 11.195 ;
      LAYER nwell ;
        RECT 77.475 10.850 79.325 13.250 ;
        RECT 80.625 10.850 82.475 13.250 ;
        RECT 8.460 6.865 10.310 9.265 ;
        RECT 12.685 6.860 21.295 9.270 ;
        RECT 23.455 6.865 25.305 9.265 ;
      LAYER pwell ;
        RECT 77.545 8.920 79.255 10.180 ;
        RECT 80.695 8.920 82.405 10.180 ;
      LAYER li1 ;
        RECT 16.565 204.145 16.965 204.495 ;
        RECT 19.665 204.345 20.170 204.645 ;
        RECT 23.365 204.195 24.120 204.580 ;
        RECT 28.165 204.395 28.760 204.700 ;
        RECT 32.365 204.200 33.115 204.595 ;
        RECT 17.295 203.540 32.215 203.800 ;
        RECT 17.295 203.065 17.695 203.540 ;
        RECT 20.445 203.065 20.845 203.540 ;
        RECT 24.220 203.070 24.620 203.540 ;
        RECT 16.245 202.725 16.645 203.065 ;
        RECT 16.165 202.265 16.645 202.725 ;
        RECT 16.895 202.265 17.695 203.065 ;
        RECT 19.395 202.725 19.795 203.065 ;
        RECT 19.315 202.265 19.795 202.725 ;
        RECT 20.045 202.265 20.845 203.065 ;
        RECT 23.170 202.815 23.570 203.070 ;
        RECT 23.085 202.270 23.570 202.815 ;
        RECT 23.820 202.270 24.620 203.070 ;
        RECT 27.560 203.075 27.960 203.540 ;
        RECT 27.560 202.275 28.360 203.075 ;
        RECT 28.610 202.275 29.015 203.075 ;
        RECT 16.165 201.545 16.565 202.265 ;
        RECT 17.015 201.545 17.340 201.620 ;
        RECT 16.165 201.345 17.340 201.545 ;
        RECT 16.165 198.955 16.565 201.345 ;
        RECT 17.015 201.295 17.340 201.345 ;
        RECT 16.815 198.955 17.615 200.755 ;
        RECT 19.315 198.955 19.715 202.265 ;
        RECT 19.965 198.955 20.765 200.755 ;
        RECT 17.265 198.555 17.615 198.955 ;
        RECT 20.415 198.555 20.765 198.955 ;
        RECT 23.085 196.855 23.485 202.270 ;
        RECT 23.735 198.950 24.535 200.750 ;
        RECT 23.740 198.555 24.535 198.950 ;
        RECT 23.740 196.855 24.530 198.555 ;
        RECT 24.165 196.470 24.530 196.855 ;
        RECT 27.565 192.925 28.365 200.855 ;
        RECT 28.615 192.930 29.015 202.275 ;
        RECT 31.815 203.070 32.215 203.540 ;
        RECT 31.815 202.270 32.615 203.070 ;
        RECT 32.865 202.270 33.265 203.070 ;
        RECT 32.870 200.855 33.265 202.270 ;
        RECT 27.565 192.600 27.970 192.925 ;
        RECT 31.815 185.030 32.615 200.850 ;
        RECT 32.865 200.055 33.265 200.855 ;
        RECT 32.870 185.030 33.265 200.055 ;
        RECT 31.815 184.730 32.215 185.030 ;
        RECT 60.500 117.560 60.670 117.645 ;
        RECT 63.220 117.560 63.390 117.645 ;
        RECT 65.940 117.560 66.110 117.645 ;
        RECT 68.660 117.560 68.830 117.645 ;
        RECT 71.380 117.560 71.550 117.645 ;
        RECT 74.100 117.560 74.270 117.645 ;
        RECT 76.820 117.560 76.990 117.645 ;
        RECT 79.540 117.560 79.710 117.645 ;
        RECT 82.260 117.560 82.430 117.645 ;
        RECT 84.980 117.560 85.150 117.645 ;
        RECT 87.700 117.560 87.870 117.645 ;
        RECT 90.420 117.560 90.590 117.645 ;
        RECT 93.140 117.560 93.310 117.645 ;
        RECT 95.860 117.560 96.030 117.645 ;
        RECT 98.580 117.560 98.750 117.645 ;
        RECT 101.300 117.560 101.470 117.645 ;
        RECT 104.020 117.560 104.190 117.645 ;
        RECT 106.740 117.560 106.910 117.645 ;
        RECT 109.460 117.560 109.630 117.645 ;
        RECT 112.180 117.560 112.350 117.645 ;
        RECT 60.500 117.040 61.960 117.560 ;
        RECT 60.500 116.350 61.420 117.040 ;
        RECT 62.130 116.870 64.480 117.560 ;
        RECT 64.650 117.040 67.400 117.560 ;
        RECT 61.590 116.350 65.020 116.870 ;
        RECT 65.190 116.350 66.860 117.040 ;
        RECT 67.570 116.870 69.920 117.560 ;
        RECT 70.090 117.040 72.840 117.560 ;
        RECT 67.030 116.350 70.460 116.870 ;
        RECT 70.630 116.350 72.300 117.040 ;
        RECT 73.010 116.870 75.360 117.560 ;
        RECT 75.530 117.040 78.280 117.560 ;
        RECT 72.470 116.350 75.900 116.870 ;
        RECT 76.070 116.350 77.740 117.040 ;
        RECT 78.450 116.870 80.800 117.560 ;
        RECT 80.970 117.040 83.720 117.560 ;
        RECT 77.910 116.350 81.340 116.870 ;
        RECT 81.510 116.350 83.180 117.040 ;
        RECT 83.890 116.870 86.240 117.560 ;
        RECT 86.410 117.040 89.160 117.560 ;
        RECT 83.350 116.350 86.780 116.870 ;
        RECT 86.950 116.350 88.620 117.040 ;
        RECT 89.330 116.870 91.680 117.560 ;
        RECT 91.850 117.040 94.600 117.560 ;
        RECT 88.790 116.350 92.220 116.870 ;
        RECT 92.390 116.350 94.060 117.040 ;
        RECT 94.770 116.870 97.120 117.560 ;
        RECT 97.290 117.040 100.040 117.560 ;
        RECT 94.230 116.350 97.660 116.870 ;
        RECT 97.830 116.350 99.500 117.040 ;
        RECT 100.210 116.870 102.560 117.560 ;
        RECT 102.730 117.040 105.480 117.560 ;
        RECT 99.670 116.350 103.100 116.870 ;
        RECT 103.270 116.350 104.940 117.040 ;
        RECT 105.650 116.870 108.000 117.560 ;
        RECT 108.170 117.040 110.920 117.560 ;
        RECT 105.110 116.350 108.540 116.870 ;
        RECT 108.710 116.350 110.380 117.040 ;
        RECT 111.090 116.870 112.350 117.560 ;
        RECT 110.550 116.350 112.350 116.870 ;
        RECT 60.500 116.180 60.670 116.350 ;
        RECT 63.220 116.180 63.390 116.350 ;
        RECT 65.940 116.180 66.110 116.350 ;
        RECT 68.660 116.180 68.830 116.350 ;
        RECT 71.380 116.180 71.550 116.350 ;
        RECT 60.500 114.970 61.960 116.180 ;
        RECT 60.500 113.590 61.440 114.970 ;
        RECT 62.130 114.800 64.480 116.180 ;
        RECT 64.650 115.430 67.400 116.180 ;
        RECT 67.570 115.490 69.920 116.180 ;
        RECT 70.090 115.660 71.550 116.180 ;
        RECT 74.100 116.180 74.270 116.350 ;
        RECT 76.820 116.180 76.990 116.350 ;
        RECT 79.540 116.180 79.710 116.350 ;
        RECT 64.650 114.970 66.880 115.430 ;
        RECT 67.570 115.260 70.460 115.490 ;
        RECT 61.610 113.590 65.000 114.800 ;
        RECT 65.170 114.510 66.880 114.970 ;
        RECT 67.050 114.970 70.460 115.260 ;
        RECT 70.630 115.290 71.550 115.660 ;
        RECT 71.975 115.525 73.325 115.695 ;
        RECT 71.975 115.460 72.305 115.525 ;
        RECT 72.960 115.395 73.325 115.525 ;
        RECT 74.100 115.490 75.360 116.180 ;
        RECT 75.530 115.660 78.280 116.180 ;
        RECT 78.450 115.740 79.710 116.180 ;
        RECT 82.260 116.180 82.430 116.350 ;
        RECT 84.980 116.180 85.150 116.350 ;
        RECT 87.700 116.180 87.870 116.350 ;
        RECT 79.880 115.920 80.810 116.100 ;
        RECT 70.630 114.970 72.290 115.290 ;
        RECT 72.460 115.005 72.790 115.350 ;
        RECT 67.050 114.510 68.830 114.970 ;
        RECT 71.380 114.960 72.290 114.970 ;
        RECT 65.170 113.590 66.110 114.510 ;
        RECT 66.280 113.620 66.830 113.790 ;
        RECT 60.500 112.990 60.670 113.590 ;
        RECT 60.930 113.160 61.390 113.330 ;
        RECT 60.500 112.660 61.050 112.990 ;
        RECT 61.220 112.895 61.390 113.160 ;
        RECT 61.560 113.065 62.210 113.415 ;
        RECT 62.380 113.160 63.050 113.330 ;
        RECT 62.380 112.895 62.550 113.160 ;
        RECT 63.220 112.990 63.390 113.590 ;
        RECT 65.940 113.440 66.110 113.590 ;
        RECT 63.560 113.160 64.230 113.330 ;
        RECT 61.220 112.665 62.550 112.895 ;
        RECT 62.720 112.660 63.890 112.990 ;
        RECT 64.060 112.895 64.230 113.160 ;
        RECT 64.400 113.065 65.050 113.415 ;
        RECT 65.220 113.160 65.680 113.330 ;
        RECT 65.220 112.895 65.390 113.160 ;
        RECT 65.940 113.110 66.490 113.440 ;
        RECT 66.660 113.295 66.830 113.620 ;
        RECT 67.010 113.520 67.380 113.860 ;
        RECT 67.560 113.620 68.490 113.800 ;
        RECT 67.560 113.295 67.730 113.620 ;
        RECT 68.660 113.440 68.830 114.510 ;
        RECT 66.660 113.125 67.730 113.295 ;
        RECT 65.940 112.990 66.110 113.110 ;
        RECT 67.085 113.020 67.415 113.125 ;
        RECT 67.900 113.110 68.830 113.440 ;
        RECT 69.050 113.140 69.340 114.800 ;
        RECT 69.510 114.475 69.970 114.800 ;
        RECT 69.510 113.375 69.680 114.475 ;
        RECT 70.140 114.445 70.710 114.800 ;
        RECT 71.380 114.795 71.550 114.960 ;
        RECT 70.880 114.460 71.550 114.795 ;
        RECT 72.960 114.775 73.130 115.395 ;
        RECT 74.100 115.225 75.900 115.490 ;
        RECT 73.300 114.970 75.900 115.225 ;
        RECT 76.070 114.970 77.740 115.660 ;
        RECT 78.450 115.490 80.470 115.740 ;
        RECT 77.910 115.410 80.470 115.490 ;
        RECT 80.640 115.595 80.810 115.920 ;
        RECT 80.990 115.820 81.360 116.160 ;
        RECT 81.540 115.920 82.090 116.090 ;
        RECT 81.540 115.595 81.710 115.920 ;
        RECT 82.260 115.740 83.720 116.180 ;
        RECT 80.640 115.425 81.710 115.595 ;
        RECT 81.880 115.430 83.720 115.740 ;
        RECT 77.910 114.970 79.710 115.410 ;
        RECT 80.955 115.320 81.285 115.425 ;
        RECT 81.880 115.410 83.200 115.430 ;
        RECT 79.880 115.150 80.785 115.240 ;
        RECT 81.585 115.150 82.090 115.230 ;
        RECT 79.880 114.970 82.090 115.150 ;
        RECT 69.850 114.275 70.020 114.280 ;
        RECT 69.850 113.565 70.470 114.275 ;
        RECT 70.640 114.090 71.160 114.260 ;
        RECT 69.510 113.205 69.970 113.375 ;
        RECT 64.060 112.665 65.390 112.895 ;
        RECT 65.560 112.660 66.110 112.990 ;
        RECT 68.660 112.970 68.830 113.110 ;
        RECT 66.280 112.850 66.785 112.930 ;
        RECT 67.585 112.850 68.490 112.940 ;
        RECT 66.280 112.670 68.490 112.850 ;
        RECT 68.660 112.690 69.630 112.970 ;
        RECT 69.800 112.820 69.970 113.205 ;
        RECT 70.140 112.990 70.470 113.395 ;
        RECT 70.640 113.390 70.810 114.090 ;
        RECT 71.380 113.890 71.550 114.460 ;
        RECT 70.980 113.560 71.550 113.890 ;
        RECT 70.640 113.220 71.160 113.390 ;
        RECT 71.380 113.360 71.550 113.560 ;
        RECT 71.720 114.450 72.370 114.725 ;
        RECT 71.720 113.780 71.930 114.450 ;
        RECT 72.540 114.445 73.130 114.775 ;
        RECT 73.300 114.440 73.930 114.770 ;
        RECT 72.100 114.275 72.400 114.280 ;
        RECT 73.300 114.275 73.470 114.440 ;
        RECT 72.100 113.995 73.470 114.275 ;
        RECT 74.100 114.305 74.270 114.970 ;
        RECT 76.820 114.795 76.990 114.970 ;
        RECT 75.045 114.605 76.395 114.775 ;
        RECT 75.045 114.475 75.410 114.605 ;
        RECT 76.065 114.540 76.395 114.605 ;
        RECT 74.100 114.270 75.070 114.305 ;
        RECT 72.100 113.950 72.370 113.995 ;
        RECT 71.720 113.530 72.370 113.780 ;
        RECT 70.640 112.820 70.810 113.220 ;
        RECT 71.380 113.190 71.990 113.360 ;
        RECT 71.380 113.050 71.550 113.190 ;
        RECT 60.500 112.050 60.670 112.660 ;
        RECT 60.930 112.305 63.050 112.490 ;
        RECT 60.500 111.800 61.130 112.050 ;
        RECT 61.300 111.855 62.250 112.135 ;
        RECT 63.220 112.065 63.390 112.660 ;
        RECT 63.560 112.305 65.680 112.490 ;
        RECT 62.760 111.800 63.850 112.065 ;
        RECT 64.360 111.855 65.310 112.135 ;
        RECT 65.940 112.070 66.110 112.660 ;
        RECT 66.370 112.240 66.830 112.410 ;
        RECT 65.940 112.050 66.490 112.070 ;
        RECT 65.480 111.800 66.490 112.050 ;
        RECT 60.500 110.105 60.670 111.800 ;
        RECT 61.260 111.630 62.625 111.685 ;
        RECT 60.950 111.515 63.050 111.630 ;
        RECT 60.950 111.460 61.390 111.515 ;
        RECT 60.950 111.295 61.120 111.460 ;
        RECT 62.495 111.380 63.050 111.515 ;
        RECT 60.950 110.595 61.120 111.100 ;
        RECT 61.320 110.935 61.540 111.290 ;
        RECT 61.710 111.105 62.305 111.345 ;
        RECT 61.320 110.765 62.605 110.935 ;
        RECT 60.950 110.425 62.070 110.595 ;
        RECT 61.900 110.235 62.070 110.425 ;
        RECT 62.240 110.405 62.605 110.765 ;
        RECT 62.775 110.235 62.945 111.170 ;
        RECT 60.500 109.735 61.170 110.105 ;
        RECT 61.350 110.015 61.680 110.215 ;
        RECT 61.900 110.065 62.945 110.235 ;
        RECT 60.500 107.920 60.670 109.735 ;
        RECT 61.350 109.555 61.650 110.015 ;
        RECT 61.900 109.895 62.160 110.065 ;
        RECT 63.220 109.895 63.390 111.800 ;
        RECT 65.940 111.740 66.490 111.800 ;
        RECT 66.660 111.975 66.830 112.240 ;
        RECT 67.000 112.145 67.650 112.495 ;
        RECT 67.820 112.240 68.490 112.410 ;
        RECT 67.820 111.975 67.990 112.240 ;
        RECT 68.660 112.070 68.830 112.690 ;
        RECT 69.800 112.650 70.810 112.820 ;
        RECT 70.980 112.670 71.550 113.050 ;
        RECT 72.160 113.020 72.370 113.530 ;
        RECT 71.720 112.670 72.370 113.020 ;
        RECT 72.540 113.625 73.120 113.815 ;
        RECT 72.540 112.670 72.740 113.625 ;
        RECT 73.300 113.525 73.470 113.995 ;
        RECT 73.640 114.050 75.070 114.270 ;
        RECT 73.640 113.695 74.270 114.050 ;
        RECT 75.240 113.855 75.410 114.475 ;
        RECT 76.820 114.460 77.490 114.795 ;
        RECT 75.580 114.085 75.910 114.430 ;
        RECT 76.820 114.370 76.990 114.460 ;
        RECT 77.660 114.445 78.230 114.800 ;
        RECT 78.400 114.475 78.860 114.800 ;
        RECT 76.080 114.040 76.990 114.370 ;
        RECT 77.210 114.090 77.730 114.260 ;
        RECT 76.820 113.890 76.990 114.040 ;
        RECT 73.300 113.445 73.930 113.525 ;
        RECT 72.960 113.170 73.930 113.445 ;
        RECT 74.100 113.350 74.270 113.695 ;
        RECT 74.440 113.520 75.070 113.850 ;
        RECT 75.240 113.525 75.830 113.855 ;
        RECT 76.000 113.530 76.650 113.805 ;
        RECT 74.900 113.355 75.070 113.520 ;
        RECT 76.100 113.355 76.270 113.360 ;
        RECT 74.100 113.000 74.730 113.350 ;
        RECT 72.960 112.775 74.730 113.000 ;
        RECT 74.900 113.075 76.270 113.355 ;
        RECT 72.960 112.670 74.270 112.775 ;
        RECT 70.140 112.545 70.470 112.650 ;
        RECT 69.000 112.375 69.970 112.480 ;
        RECT 70.705 112.375 71.050 112.480 ;
        RECT 69.000 112.205 71.050 112.375 ;
        RECT 66.660 111.745 67.990 111.975 ;
        RECT 68.160 112.035 68.830 112.070 ;
        RECT 71.380 112.070 71.550 112.670 ;
        RECT 71.810 112.240 72.270 112.410 ;
        RECT 71.380 112.035 71.930 112.070 ;
        RECT 68.160 111.865 70.010 112.035 ;
        RECT 70.465 111.865 71.930 112.035 ;
        RECT 68.160 111.740 68.830 111.865 ;
        RECT 63.985 111.630 65.350 111.685 ;
        RECT 63.560 111.515 65.660 111.630 ;
        RECT 63.560 111.380 64.115 111.515 ;
        RECT 65.220 111.460 65.660 111.515 ;
        RECT 63.665 110.235 63.835 111.170 ;
        RECT 64.305 111.105 64.900 111.345 ;
        RECT 65.490 111.295 65.660 111.460 ;
        RECT 65.070 110.935 65.290 111.290 ;
        RECT 65.940 111.130 66.110 111.740 ;
        RECT 66.370 111.385 68.490 111.570 ;
        RECT 64.005 110.765 65.290 110.935 ;
        RECT 64.005 110.405 64.370 110.765 ;
        RECT 65.490 110.595 65.660 111.100 ;
        RECT 64.540 110.425 65.660 110.595 ;
        RECT 65.940 110.880 66.570 111.130 ;
        RECT 66.740 110.935 67.690 111.215 ;
        RECT 68.660 111.145 68.830 111.740 ;
        RECT 71.380 111.740 71.930 111.865 ;
        RECT 72.100 111.975 72.270 112.240 ;
        RECT 72.440 112.145 73.090 112.495 ;
        RECT 73.260 112.240 73.930 112.410 ;
        RECT 73.260 111.975 73.430 112.240 ;
        RECT 74.100 112.080 74.270 112.670 ;
        RECT 74.900 112.605 75.070 113.075 ;
        RECT 76.000 113.030 76.270 113.075 ;
        RECT 75.290 112.895 75.460 112.900 ;
        RECT 75.250 112.705 75.830 112.895 ;
        RECT 76.440 112.860 76.650 113.530 ;
        RECT 74.440 112.525 75.070 112.605 ;
        RECT 74.440 112.250 75.410 112.525 ;
        RECT 74.100 112.070 75.410 112.080 ;
        RECT 72.100 111.745 73.430 111.975 ;
        RECT 73.600 111.750 75.410 112.070 ;
        RECT 75.630 111.750 75.830 112.705 ;
        RECT 76.000 112.610 76.650 112.860 ;
        RECT 76.820 113.560 77.390 113.890 ;
        RECT 76.820 113.050 76.990 113.560 ;
        RECT 77.560 113.390 77.730 114.090 ;
        RECT 77.900 113.565 78.520 114.275 ;
        RECT 77.210 113.220 77.730 113.390 ;
        RECT 76.820 112.670 77.390 113.050 ;
        RECT 77.560 112.820 77.730 113.220 ;
        RECT 77.900 112.990 78.230 113.395 ;
        RECT 78.690 113.375 78.860 114.475 ;
        RECT 78.400 113.205 78.860 113.375 ;
        RECT 78.400 112.820 78.570 113.205 ;
        RECT 79.030 113.140 79.320 114.800 ;
        RECT 79.540 114.360 79.710 114.970 ;
        RECT 79.880 114.540 80.810 114.720 ;
        RECT 79.540 114.030 80.470 114.360 ;
        RECT 80.640 114.215 80.810 114.540 ;
        RECT 80.990 114.440 81.360 114.780 ;
        RECT 81.540 114.540 82.090 114.710 ;
        RECT 81.540 114.215 81.710 114.540 ;
        RECT 82.260 114.510 83.200 115.410 ;
        RECT 83.890 115.260 85.585 116.180 ;
        RECT 83.370 114.510 85.585 115.260 ;
        RECT 87.155 115.740 87.870 116.180 ;
        RECT 88.040 115.920 88.590 116.090 ;
        RECT 87.155 115.410 88.250 115.740 ;
        RECT 88.420 115.595 88.590 115.920 ;
        RECT 88.770 115.820 89.140 116.160 ;
        RECT 89.320 115.920 90.250 116.100 ;
        RECT 89.320 115.595 89.490 115.920 ;
        RECT 90.420 115.740 90.590 116.350 ;
        RECT 93.140 116.180 93.310 116.350 ;
        RECT 95.860 116.180 96.030 116.350 ;
        RECT 98.580 116.180 98.750 116.350 ;
        RECT 101.300 116.180 101.470 116.350 ;
        RECT 90.760 115.920 91.690 116.100 ;
        RECT 88.420 115.425 89.490 115.595 ;
        RECT 87.155 114.595 87.870 115.410 ;
        RECT 88.845 115.320 89.175 115.425 ;
        RECT 89.660 115.410 91.350 115.740 ;
        RECT 91.520 115.595 91.690 115.920 ;
        RECT 91.870 115.820 92.240 116.160 ;
        RECT 92.420 115.920 92.970 116.090 ;
        RECT 92.420 115.595 92.590 115.920 ;
        RECT 93.140 115.740 93.855 116.180 ;
        RECT 91.520 115.425 92.590 115.595 ;
        RECT 88.040 115.150 88.545 115.230 ;
        RECT 89.345 115.150 90.250 115.240 ;
        RECT 88.040 114.970 90.250 115.150 ;
        RECT 82.260 114.360 82.430 114.510 ;
        RECT 80.640 114.045 81.710 114.215 ;
        RECT 79.540 112.990 79.710 114.030 ;
        RECT 80.955 113.940 81.285 114.045 ;
        RECT 81.880 114.030 82.430 114.360 ;
        RECT 79.880 113.770 80.785 113.860 ;
        RECT 81.585 113.770 82.090 113.850 ;
        RECT 79.880 113.590 82.090 113.770 ;
        RECT 82.260 113.450 82.430 114.030 ;
        RECT 82.690 113.620 83.150 113.790 ;
        RECT 79.880 113.160 80.550 113.330 ;
        RECT 79.540 112.970 80.210 112.990 ;
        RECT 76.000 112.100 76.210 112.610 ;
        RECT 76.820 112.440 76.990 112.670 ;
        RECT 77.560 112.650 78.570 112.820 ;
        RECT 78.740 112.690 80.210 112.970 ;
        RECT 79.540 112.660 80.210 112.690 ;
        RECT 80.380 112.895 80.550 113.160 ;
        RECT 80.720 113.065 81.370 113.415 ;
        RECT 81.540 113.160 82.000 113.330 ;
        RECT 81.540 112.895 81.710 113.160 ;
        RECT 82.260 113.120 82.810 113.450 ;
        RECT 82.980 113.355 83.150 113.620 ;
        RECT 83.320 113.525 83.970 113.875 ;
        RECT 84.140 113.620 84.810 113.790 ;
        RECT 84.140 113.355 84.310 113.620 ;
        RECT 84.980 113.450 85.585 114.510 ;
        RECT 86.325 114.370 87.870 114.595 ;
        RECT 88.130 114.540 88.590 114.710 ;
        RECT 86.325 114.255 88.250 114.370 ;
        RECT 82.980 113.125 84.310 113.355 ;
        RECT 84.480 113.120 85.585 113.450 ;
        RECT 82.260 112.990 82.430 113.120 ;
        RECT 80.380 112.665 81.710 112.895 ;
        RECT 81.880 112.660 82.430 112.990 ;
        RECT 82.690 112.765 84.810 112.950 ;
        RECT 84.980 112.775 85.585 113.120 ;
        RECT 87.155 114.040 88.250 114.255 ;
        RECT 88.420 114.275 88.590 114.540 ;
        RECT 88.760 114.445 89.410 114.795 ;
        RECT 89.580 114.540 90.250 114.710 ;
        RECT 89.580 114.275 89.750 114.540 ;
        RECT 90.420 114.370 90.590 115.410 ;
        RECT 91.835 115.320 92.165 115.425 ;
        RECT 92.760 115.410 93.855 115.740 ;
        RECT 90.760 115.150 91.665 115.240 ;
        RECT 92.465 115.150 92.970 115.230 ;
        RECT 90.760 114.970 92.970 115.150 ;
        RECT 90.760 114.540 91.430 114.710 ;
        RECT 88.420 114.045 89.750 114.275 ;
        RECT 89.920 114.040 91.090 114.370 ;
        RECT 91.260 114.275 91.430 114.540 ;
        RECT 91.600 114.445 92.250 114.795 ;
        RECT 92.420 114.540 92.880 114.710 ;
        RECT 93.140 114.595 93.855 115.410 ;
        RECT 95.425 115.490 97.120 116.180 ;
        RECT 97.290 115.660 100.040 116.180 ;
        RECT 95.425 114.970 97.660 115.490 ;
        RECT 97.830 115.430 100.040 115.660 ;
        RECT 100.210 115.740 101.470 116.180 ;
        RECT 101.640 115.920 102.570 116.100 ;
        RECT 97.830 114.970 99.520 115.430 ;
        RECT 100.210 115.410 102.230 115.740 ;
        RECT 102.400 115.595 102.570 115.920 ;
        RECT 102.750 115.820 103.120 116.160 ;
        RECT 103.300 115.920 103.850 116.090 ;
        RECT 103.300 115.595 103.470 115.920 ;
        RECT 104.020 115.740 104.190 116.350 ;
        RECT 102.400 115.425 103.470 115.595 ;
        RECT 100.210 115.260 101.470 115.410 ;
        RECT 102.715 115.320 103.045 115.425 ;
        RECT 103.640 115.410 104.190 115.740 ;
        RECT 92.420 114.275 92.590 114.540 ;
        RECT 93.140 114.370 94.685 114.595 ;
        RECT 91.260 114.045 92.590 114.275 ;
        RECT 92.760 114.255 94.685 114.370 ;
        RECT 92.760 114.040 93.855 114.255 ;
        RECT 87.155 113.430 87.870 114.040 ;
        RECT 88.130 113.685 90.250 113.870 ;
        RECT 87.155 113.180 88.330 113.430 ;
        RECT 88.500 113.235 89.450 113.515 ;
        RECT 90.420 113.445 90.590 114.040 ;
        RECT 90.760 113.685 92.880 113.870 ;
        RECT 89.960 113.180 91.050 113.445 ;
        RECT 91.560 113.235 92.510 113.515 ;
        RECT 93.140 113.430 93.855 114.040 ;
        RECT 92.680 113.180 93.855 113.430 ;
        RECT 77.900 112.545 78.230 112.650 ;
        RECT 76.380 112.270 76.990 112.440 ;
        RECT 76.000 111.750 76.650 112.100 ;
        RECT 76.820 112.035 76.990 112.270 ;
        RECT 77.320 112.375 77.665 112.480 ;
        RECT 78.400 112.375 79.370 112.480 ;
        RECT 77.320 112.205 79.370 112.375 ;
        RECT 79.540 112.065 79.710 112.660 ;
        RECT 82.260 112.510 82.430 112.660 ;
        RECT 79.880 112.305 82.000 112.490 ;
        RECT 82.260 112.260 82.890 112.510 ;
        RECT 83.060 112.315 84.010 112.595 ;
        RECT 84.980 112.525 86.835 112.775 ;
        RECT 84.520 112.425 86.835 112.525 ;
        RECT 84.520 112.260 85.585 112.425 ;
        RECT 79.540 112.035 80.170 112.065 ;
        RECT 76.820 111.865 77.905 112.035 ;
        RECT 78.360 111.865 80.170 112.035 ;
        RECT 73.600 111.740 74.270 111.750 ;
        RECT 69.000 111.320 69.930 111.500 ;
        RECT 68.200 111.140 68.830 111.145 ;
        RECT 68.200 110.880 69.590 111.140 ;
        RECT 64.540 110.235 64.710 110.425 ;
        RECT 63.665 110.065 64.710 110.235 ;
        RECT 64.450 109.895 64.710 110.065 ;
        RECT 64.930 110.015 65.260 110.215 ;
        RECT 65.940 110.105 66.110 110.880 ;
        RECT 68.660 110.810 69.590 110.880 ;
        RECT 69.760 110.995 69.930 111.320 ;
        RECT 70.110 111.220 70.480 111.560 ;
        RECT 70.660 111.320 71.210 111.490 ;
        RECT 70.660 110.995 70.830 111.320 ;
        RECT 71.380 111.140 71.550 111.740 ;
        RECT 71.810 111.385 73.930 111.570 ;
        RECT 69.760 110.825 70.830 110.995 ;
        RECT 71.000 111.130 71.550 111.140 ;
        RECT 71.000 110.880 72.010 111.130 ;
        RECT 72.180 110.935 73.130 111.215 ;
        RECT 74.100 111.145 74.270 111.740 ;
        RECT 76.820 111.580 76.990 111.865 ;
        RECT 79.540 111.800 80.170 111.865 ;
        RECT 80.680 111.855 81.630 112.135 ;
        RECT 82.260 112.050 82.430 112.260 ;
        RECT 83.020 112.090 84.385 112.145 ;
        RECT 81.800 111.800 82.430 112.050 ;
        RECT 79.540 111.580 79.710 111.800 ;
        RECT 80.305 111.630 81.670 111.685 ;
        RECT 73.640 110.880 74.270 111.145 ;
        RECT 66.700 110.710 68.065 110.765 ;
        RECT 66.390 110.595 68.490 110.710 ;
        RECT 66.390 110.540 66.830 110.595 ;
        RECT 66.390 110.375 66.560 110.540 ;
        RECT 67.935 110.460 68.490 110.595 ;
        RECT 61.830 109.725 62.160 109.895 ;
        RECT 62.420 109.725 64.190 109.895 ;
        RECT 64.450 109.725 64.780 109.895 ;
        RECT 60.950 109.385 63.050 109.555 ;
        RECT 60.950 109.150 61.120 109.385 ;
        RECT 62.720 109.305 63.050 109.385 ;
        RECT 61.830 109.025 62.550 109.215 ;
        RECT 60.950 108.365 61.120 108.980 ;
        RECT 61.290 108.855 61.620 109.000 ;
        RECT 61.290 108.535 62.580 108.855 ;
        RECT 62.750 108.365 62.920 109.080 ;
        RECT 60.950 108.195 62.920 108.365 ;
        RECT 60.500 107.710 61.200 107.920 ;
        RECT 60.500 106.950 60.670 107.710 ;
        RECT 61.580 107.490 61.910 108.195 ;
        RECT 62.115 107.470 62.490 108.025 ;
        RECT 63.220 108.015 63.390 109.725 ;
        RECT 64.960 109.555 65.260 110.015 ;
        RECT 65.440 109.735 66.110 110.105 ;
        RECT 63.560 109.385 65.660 109.555 ;
        RECT 63.560 109.305 63.890 109.385 ;
        RECT 63.690 108.365 63.860 109.080 ;
        RECT 64.060 109.025 64.780 109.215 ;
        RECT 65.490 109.150 65.660 109.385 ;
        RECT 65.940 109.185 66.110 109.735 ;
        RECT 66.390 109.675 66.560 110.180 ;
        RECT 66.760 110.015 66.980 110.370 ;
        RECT 67.150 110.185 67.745 110.425 ;
        RECT 66.760 109.845 68.045 110.015 ;
        RECT 66.390 109.505 67.510 109.675 ;
        RECT 67.340 109.315 67.510 109.505 ;
        RECT 67.680 109.485 68.045 109.845 ;
        RECT 68.215 109.315 68.385 110.250 ;
        RECT 64.990 108.855 65.320 109.000 ;
        RECT 64.030 108.535 65.320 108.855 ;
        RECT 65.490 108.365 65.660 108.980 ;
        RECT 63.690 108.195 65.660 108.365 ;
        RECT 65.940 108.815 66.610 109.185 ;
        RECT 66.790 109.095 67.120 109.295 ;
        RECT 67.340 109.145 68.385 109.315 ;
        RECT 68.660 110.200 68.830 110.810 ;
        RECT 70.075 110.720 70.405 110.825 ;
        RECT 71.000 110.810 71.550 110.880 ;
        RECT 69.000 110.550 69.905 110.640 ;
        RECT 70.705 110.550 71.210 110.630 ;
        RECT 69.000 110.370 71.210 110.550 ;
        RECT 71.380 110.200 71.550 110.810 ;
        RECT 72.140 110.710 73.505 110.765 ;
        RECT 71.830 110.595 73.930 110.710 ;
        RECT 71.830 110.540 72.270 110.595 ;
        RECT 71.830 110.375 72.000 110.540 ;
        RECT 73.375 110.460 73.930 110.595 ;
        RECT 62.720 107.700 63.890 108.015 ;
        RECT 60.885 107.320 61.410 107.450 ;
        RECT 62.115 107.320 63.050 107.470 ;
        RECT 60.885 107.130 63.050 107.320 ;
        RECT 60.885 107.120 61.910 107.130 ;
        RECT 60.500 106.780 61.280 106.950 ;
        RECT 60.500 106.110 60.670 106.780 ;
        RECT 60.890 106.455 61.410 106.610 ;
        RECT 61.580 106.570 61.910 107.120 ;
        RECT 63.220 106.960 63.390 107.700 ;
        RECT 64.120 107.470 64.495 108.025 ;
        RECT 64.700 107.490 65.030 108.195 ;
        RECT 65.940 107.920 66.110 108.815 ;
        RECT 66.790 108.635 67.090 109.095 ;
        RECT 67.340 108.975 67.600 109.145 ;
        RECT 68.660 108.975 69.920 110.200 ;
        RECT 67.270 108.805 67.600 108.975 ;
        RECT 67.860 108.805 69.920 108.975 ;
        RECT 66.390 108.465 68.490 108.635 ;
        RECT 66.390 108.230 66.560 108.465 ;
        RECT 68.160 108.385 68.490 108.465 ;
        RECT 68.660 108.380 69.920 108.805 ;
        RECT 70.090 109.185 71.550 110.200 ;
        RECT 71.830 109.675 72.000 110.180 ;
        RECT 72.200 110.015 72.420 110.370 ;
        RECT 72.590 110.185 73.185 110.425 ;
        RECT 72.200 109.845 73.485 110.015 ;
        RECT 71.830 109.505 72.950 109.675 ;
        RECT 72.780 109.315 72.950 109.505 ;
        RECT 73.120 109.485 73.485 109.845 ;
        RECT 73.655 109.315 73.825 110.250 ;
        RECT 70.090 108.815 72.050 109.185 ;
        RECT 72.230 109.095 72.560 109.295 ;
        RECT 72.780 109.145 73.825 109.315 ;
        RECT 74.100 110.215 74.270 110.880 ;
        RECT 74.490 110.385 74.780 111.580 ;
        RECT 74.950 111.230 75.410 111.560 ;
        RECT 75.580 111.230 75.910 111.580 ;
        RECT 76.080 111.305 76.600 111.560 ;
        RECT 74.950 110.565 75.120 111.230 ;
        RECT 75.290 110.835 75.910 111.060 ;
        RECT 74.950 110.395 75.410 110.565 ;
        RECT 74.100 109.935 75.070 110.215 ;
        RECT 75.240 110.065 75.410 110.395 ;
        RECT 75.580 110.235 75.910 110.835 ;
        RECT 76.080 110.635 76.250 111.305 ;
        RECT 76.820 111.135 77.535 111.580 ;
        RECT 76.420 110.805 77.535 111.135 ;
        RECT 76.080 110.465 76.600 110.635 ;
        RECT 76.080 110.065 76.250 110.465 ;
        RECT 76.820 110.295 77.535 110.805 ;
        RECT 74.100 109.280 74.270 109.935 ;
        RECT 75.240 109.895 76.250 110.065 ;
        RECT 76.420 109.995 77.535 110.295 ;
        RECT 76.420 109.915 78.365 109.995 ;
        RECT 75.580 109.790 75.910 109.895 ;
        RECT 74.440 109.620 75.410 109.725 ;
        RECT 76.145 109.620 76.490 109.725 ;
        RECT 74.440 109.450 76.490 109.620 ;
        RECT 76.820 109.655 78.365 109.915 ;
        RECT 79.105 109.895 79.710 111.580 ;
        RECT 79.880 111.515 81.980 111.630 ;
        RECT 79.880 111.380 80.435 111.515 ;
        RECT 81.540 111.460 81.980 111.515 ;
        RECT 79.985 110.235 80.155 111.170 ;
        RECT 80.625 111.105 81.220 111.345 ;
        RECT 81.810 111.295 81.980 111.460 ;
        RECT 81.390 110.935 81.610 111.290 ;
        RECT 80.325 110.765 81.610 110.935 ;
        RECT 80.325 110.405 80.690 110.765 ;
        RECT 81.810 110.595 81.980 111.100 ;
        RECT 80.860 110.425 81.980 110.595 ;
        RECT 82.260 110.565 82.430 111.800 ;
        RECT 82.710 111.975 84.810 112.090 ;
        RECT 82.710 111.920 83.150 111.975 ;
        RECT 82.710 111.755 82.880 111.920 ;
        RECT 84.255 111.840 84.810 111.975 ;
        RECT 82.710 111.055 82.880 111.560 ;
        RECT 83.080 111.395 83.300 111.750 ;
        RECT 83.470 111.565 84.065 111.805 ;
        RECT 83.080 111.225 84.365 111.395 ;
        RECT 82.710 110.885 83.830 111.055 ;
        RECT 83.660 110.695 83.830 110.885 ;
        RECT 84.000 110.865 84.365 111.225 ;
        RECT 84.535 110.695 84.705 111.630 ;
        RECT 80.860 110.235 81.030 110.425 ;
        RECT 79.985 110.065 81.030 110.235 ;
        RECT 80.770 109.895 81.030 110.065 ;
        RECT 81.250 110.015 81.580 110.215 ;
        RECT 82.260 110.195 82.930 110.565 ;
        RECT 83.110 110.475 83.440 110.675 ;
        RECT 83.660 110.525 84.705 110.695 ;
        RECT 84.980 110.835 85.585 112.260 ;
        RECT 87.155 111.485 87.870 113.180 ;
        RECT 88.460 113.010 89.825 113.065 ;
        RECT 88.150 112.895 90.250 113.010 ;
        RECT 88.150 112.840 88.590 112.895 ;
        RECT 88.150 112.675 88.320 112.840 ;
        RECT 89.695 112.760 90.250 112.895 ;
        RECT 88.150 111.975 88.320 112.480 ;
        RECT 88.520 112.315 88.740 112.670 ;
        RECT 88.910 112.485 89.505 112.725 ;
        RECT 88.520 112.145 89.805 112.315 ;
        RECT 88.150 111.805 89.270 111.975 ;
        RECT 89.100 111.615 89.270 111.805 ;
        RECT 89.440 111.785 89.805 112.145 ;
        RECT 89.975 111.615 90.145 112.550 ;
        RECT 87.155 111.115 88.370 111.485 ;
        RECT 88.550 111.395 88.880 111.595 ;
        RECT 89.100 111.445 90.145 111.615 ;
        RECT 87.155 110.835 87.870 111.115 ;
        RECT 88.550 110.935 88.850 111.395 ;
        RECT 89.100 111.275 89.360 111.445 ;
        RECT 90.420 111.275 90.590 113.180 ;
        RECT 91.185 113.010 92.550 113.065 ;
        RECT 90.760 112.895 92.860 113.010 ;
        RECT 90.760 112.760 91.315 112.895 ;
        RECT 92.420 112.840 92.860 112.895 ;
        RECT 90.865 111.615 91.035 112.550 ;
        RECT 91.505 112.485 92.100 112.725 ;
        RECT 92.690 112.675 92.860 112.840 ;
        RECT 92.270 112.315 92.490 112.670 ;
        RECT 91.205 112.145 92.490 112.315 ;
        RECT 91.205 111.785 91.570 112.145 ;
        RECT 92.690 111.975 92.860 112.480 ;
        RECT 91.740 111.805 92.860 111.975 ;
        RECT 91.740 111.615 91.910 111.805 ;
        RECT 90.865 111.445 91.910 111.615 ;
        RECT 91.650 111.275 91.910 111.445 ;
        RECT 92.130 111.395 92.460 111.595 ;
        RECT 93.140 111.485 93.855 113.180 ;
        RECT 95.425 112.970 96.030 114.970 ;
        RECT 96.250 113.140 96.540 114.800 ;
        RECT 96.710 114.475 97.170 114.800 ;
        RECT 96.710 113.375 96.880 114.475 ;
        RECT 97.340 114.445 97.910 114.800 ;
        RECT 98.580 114.795 99.520 114.970 ;
        RECT 98.080 114.510 99.520 114.795 ;
        RECT 99.690 114.510 101.470 115.260 ;
        RECT 101.640 115.150 102.545 115.240 ;
        RECT 103.345 115.150 103.850 115.230 ;
        RECT 101.640 114.970 103.850 115.150 ;
        RECT 104.020 114.820 104.190 115.410 ;
        RECT 106.740 116.180 106.910 116.350 ;
        RECT 109.460 116.180 109.630 116.350 ;
        RECT 112.180 116.180 112.350 116.350 ;
        RECT 104.360 115.000 104.910 115.170 ;
        RECT 101.640 114.540 102.570 114.720 ;
        RECT 98.080 114.460 98.750 114.510 ;
        RECT 97.050 114.275 97.220 114.280 ;
        RECT 97.050 113.565 97.670 114.275 ;
        RECT 97.840 114.090 98.360 114.260 ;
        RECT 96.710 113.205 97.170 113.375 ;
        RECT 95.425 112.775 96.830 112.970 ;
        RECT 94.175 112.690 96.830 112.775 ;
        RECT 97.000 112.820 97.170 113.205 ;
        RECT 97.340 112.990 97.670 113.395 ;
        RECT 97.840 113.390 98.010 114.090 ;
        RECT 98.580 113.910 98.750 114.460 ;
        RECT 101.300 114.360 101.470 114.510 ;
        RECT 99.010 114.080 99.470 114.250 ;
        RECT 98.580 113.890 99.130 113.910 ;
        RECT 98.180 113.580 99.130 113.890 ;
        RECT 99.300 113.815 99.470 114.080 ;
        RECT 99.640 113.985 100.290 114.335 ;
        RECT 100.460 114.080 101.130 114.250 ;
        RECT 100.460 113.815 100.630 114.080 ;
        RECT 101.300 114.030 102.230 114.360 ;
        RECT 102.400 114.215 102.570 114.540 ;
        RECT 102.750 114.440 103.120 114.780 ;
        RECT 103.300 114.540 103.850 114.710 ;
        RECT 103.300 114.215 103.470 114.540 ;
        RECT 104.020 114.490 104.570 114.820 ;
        RECT 104.740 114.675 104.910 115.000 ;
        RECT 105.090 114.900 105.460 115.240 ;
        RECT 105.640 115.000 106.570 115.180 ;
        RECT 105.640 114.675 105.810 115.000 ;
        RECT 106.740 114.820 108.000 116.180 ;
        RECT 108.170 114.970 110.175 116.180 ;
        RECT 104.740 114.505 105.810 114.675 ;
        RECT 105.980 114.800 108.000 114.820 ;
        RECT 104.020 114.360 104.190 114.490 ;
        RECT 105.165 114.400 105.495 114.505 ;
        RECT 105.980 114.490 108.520 114.800 ;
        RECT 102.400 114.045 103.470 114.215 ;
        RECT 101.300 113.910 101.470 114.030 ;
        RECT 102.715 113.940 103.045 114.045 ;
        RECT 103.640 114.030 104.190 114.360 ;
        RECT 104.360 114.230 104.865 114.310 ;
        RECT 105.665 114.230 106.570 114.320 ;
        RECT 104.360 114.050 106.570 114.230 ;
        RECT 99.300 113.585 100.630 113.815 ;
        RECT 100.800 113.580 101.470 113.910 ;
        RECT 101.640 113.770 102.545 113.860 ;
        RECT 103.345 113.770 103.850 113.850 ;
        RECT 101.640 113.590 103.850 113.770 ;
        RECT 98.180 113.560 98.750 113.580 ;
        RECT 97.840 113.220 98.360 113.390 ;
        RECT 97.840 112.820 98.010 113.220 ;
        RECT 98.580 113.050 98.750 113.560 ;
        RECT 99.010 113.225 101.130 113.410 ;
        RECT 94.175 112.425 96.030 112.690 ;
        RECT 97.000 112.650 98.010 112.820 ;
        RECT 98.180 112.970 98.750 113.050 ;
        RECT 98.180 112.720 99.210 112.970 ;
        RECT 99.380 112.775 100.330 113.055 ;
        RECT 101.300 112.990 101.470 113.580 ;
        RECT 104.020 113.450 104.190 114.030 ;
        RECT 104.450 113.620 104.910 113.790 ;
        RECT 101.640 113.160 102.310 113.330 ;
        RECT 101.300 112.985 101.970 112.990 ;
        RECT 100.840 112.720 101.970 112.985 ;
        RECT 98.180 112.670 98.750 112.720 ;
        RECT 97.340 112.545 97.670 112.650 ;
        RECT 89.030 111.105 89.360 111.275 ;
        RECT 89.620 111.105 91.390 111.275 ;
        RECT 91.650 111.105 91.980 111.275 ;
        RECT 84.980 110.660 85.150 110.835 ;
        RECT 87.700 110.660 87.870 110.835 ;
        RECT 82.260 110.105 82.430 110.195 ;
        RECT 79.105 109.725 80.510 109.895 ;
        RECT 80.770 109.725 81.100 109.895 ;
        RECT 76.820 109.280 77.535 109.655 ;
        RECT 70.090 108.550 71.550 108.815 ;
        RECT 72.230 108.635 72.530 109.095 ;
        RECT 72.780 108.975 73.040 109.145 ;
        RECT 74.100 108.990 75.475 109.280 ;
        RECT 75.990 108.990 77.535 109.280 ;
        RECT 74.100 108.975 74.270 108.990 ;
        RECT 72.710 108.805 73.040 108.975 ;
        RECT 73.300 108.820 74.270 108.975 ;
        RECT 76.820 108.820 77.535 108.990 ;
        RECT 73.300 108.805 74.705 108.820 ;
        RECT 67.270 108.105 67.990 108.295 ;
        RECT 65.410 107.710 66.110 107.920 ;
        RECT 63.560 107.320 64.495 107.470 ;
        RECT 65.200 107.320 65.725 107.450 ;
        RECT 63.560 107.130 65.725 107.320 ;
        RECT 64.700 107.120 65.725 107.130 ;
        RECT 62.210 106.790 64.400 106.960 ;
        RECT 60.890 106.400 61.450 106.455 ;
        RECT 62.080 106.445 63.005 106.620 ;
        RECT 62.030 106.400 63.005 106.445 ;
        RECT 60.890 106.290 63.005 106.400 ;
        RECT 60.890 106.280 62.160 106.290 ;
        RECT 61.325 106.230 62.160 106.280 ;
        RECT 63.220 106.120 63.390 106.790 ;
        RECT 63.605 106.445 64.530 106.620 ;
        RECT 64.700 106.570 65.030 107.120 ;
        RECT 65.940 107.000 66.110 107.710 ;
        RECT 66.390 107.445 66.560 108.060 ;
        RECT 66.730 107.935 67.060 108.080 ;
        RECT 66.730 107.615 68.020 107.935 ;
        RECT 68.190 107.445 68.360 108.160 ;
        RECT 66.390 107.275 68.360 107.445 ;
        RECT 65.940 106.950 66.640 107.000 ;
        RECT 65.330 106.790 66.640 106.950 ;
        RECT 65.330 106.780 66.110 106.790 ;
        RECT 65.200 106.455 65.720 106.610 ;
        RECT 63.605 106.400 64.580 106.445 ;
        RECT 65.160 106.400 65.720 106.455 ;
        RECT 63.605 106.290 65.720 106.400 ;
        RECT 64.450 106.280 65.720 106.290 ;
        RECT 64.450 106.230 65.285 106.280 ;
        RECT 60.500 105.940 61.185 106.110 ;
        RECT 62.305 105.950 64.305 106.120 ;
        RECT 65.940 106.110 66.110 106.780 ;
        RECT 67.020 106.570 67.350 107.275 ;
        RECT 67.555 106.550 67.930 107.105 ;
        RECT 68.660 107.095 70.440 108.380 ;
        RECT 68.160 106.780 70.440 107.095 ;
        RECT 68.660 106.690 70.440 106.780 ;
        RECT 70.610 107.000 71.550 108.550 ;
        RECT 71.830 108.465 73.930 108.635 ;
        RECT 71.830 108.230 72.000 108.465 ;
        RECT 73.600 108.385 73.930 108.465 ;
        RECT 72.710 108.105 73.430 108.295 ;
        RECT 71.830 107.445 72.000 108.060 ;
        RECT 72.170 107.935 72.500 108.080 ;
        RECT 72.170 107.615 73.460 107.935 ;
        RECT 73.630 107.445 73.800 108.160 ;
        RECT 71.830 107.275 73.800 107.445 ;
        RECT 70.610 106.790 72.080 107.000 ;
        RECT 70.610 106.690 71.550 106.790 ;
        RECT 66.325 106.400 66.850 106.530 ;
        RECT 67.555 106.400 68.490 106.550 ;
        RECT 66.325 106.210 68.490 106.400 ;
        RECT 68.660 106.500 68.830 106.690 ;
        RECT 66.325 106.200 67.350 106.210 ;
        RECT 65.425 106.030 66.110 106.110 ;
        RECT 60.500 104.680 60.670 105.940 ;
        RECT 63.220 105.600 63.390 105.950 ;
        RECT 65.425 105.940 66.720 106.030 ;
        RECT 65.940 105.860 66.720 105.940 ;
        RECT 65.940 105.600 66.110 105.860 ;
        RECT 63.220 104.680 64.480 105.600 ;
        RECT 64.650 105.190 66.110 105.600 ;
        RECT 66.330 105.535 66.850 105.690 ;
        RECT 67.020 105.650 67.350 106.200 ;
        RECT 68.660 106.170 69.680 106.500 ;
        RECT 68.660 106.040 68.830 106.170 ;
        RECT 67.650 105.870 68.830 106.040 ;
        RECT 69.850 106.155 70.410 106.485 ;
        RECT 70.580 106.170 71.210 106.500 ;
        RECT 66.330 105.480 66.890 105.535 ;
        RECT 67.520 105.525 68.445 105.700 ;
        RECT 67.470 105.480 68.445 105.525 ;
        RECT 66.330 105.370 68.445 105.480 ;
        RECT 66.330 105.360 67.600 105.370 ;
        RECT 66.765 105.310 67.600 105.360 ;
        RECT 68.660 105.200 68.830 105.870 ;
        RECT 64.650 105.020 66.625 105.190 ;
        RECT 67.745 105.030 68.830 105.200 ;
        RECT 64.650 104.850 66.110 105.020 ;
        RECT 65.170 104.680 66.110 104.850 ;
        RECT 68.660 104.695 68.830 105.030 ;
        RECT 69.000 105.780 69.680 106.000 ;
        RECT 69.000 105.080 69.170 105.780 ;
        RECT 69.340 105.310 69.680 105.610 ;
        RECT 69.000 104.890 69.330 105.080 ;
        RECT 68.660 104.680 69.290 104.695 ;
        RECT 60.500 104.390 61.395 104.680 ;
        RECT 62.055 104.390 65.000 104.680 ;
        RECT 60.500 104.220 60.670 104.390 ;
        RECT 63.220 104.220 65.000 104.390 ;
        RECT 60.500 102.635 61.215 104.220 ;
        RECT 62.785 103.930 65.000 104.220 ;
        RECT 65.170 104.390 66.835 104.680 ;
        RECT 67.495 104.390 69.290 104.680 ;
        RECT 65.170 103.930 66.110 104.390 ;
        RECT 62.785 103.655 63.390 103.930 ;
        RECT 62.785 103.485 63.850 103.655 ;
        RECT 62.785 102.815 63.390 103.485 ;
        RECT 64.020 103.330 65.370 103.760 ;
        RECT 65.940 103.735 66.110 103.930 ;
        RECT 65.540 103.405 66.110 103.735 ;
        RECT 64.020 103.315 64.190 103.330 ;
        RECT 63.560 102.985 64.190 103.315 ;
        RECT 65.200 103.235 65.370 103.330 ;
        RECT 65.940 103.295 66.110 103.405 ;
        RECT 68.660 104.365 69.290 104.390 ;
        RECT 68.660 103.790 68.830 104.365 ;
        RECT 69.500 104.195 69.680 105.310 ;
        RECT 69.850 105.005 70.020 106.155 ;
        RECT 70.190 105.185 70.390 105.985 ;
        RECT 70.580 105.640 70.750 106.170 ;
        RECT 71.380 106.030 71.550 106.690 ;
        RECT 72.460 106.570 72.790 107.275 ;
        RECT 72.995 106.550 73.370 107.105 ;
        RECT 74.100 107.095 74.705 108.805 ;
        RECT 76.275 107.235 77.535 108.820 ;
        RECT 79.105 108.175 79.710 109.725 ;
        RECT 81.280 109.555 81.580 110.015 ;
        RECT 81.760 109.735 82.430 110.105 ;
        RECT 83.110 110.015 83.410 110.475 ;
        RECT 83.660 110.355 83.920 110.525 ;
        RECT 84.980 110.355 86.240 110.660 ;
        RECT 83.590 110.185 83.920 110.355 ;
        RECT 84.180 110.185 86.240 110.355 ;
        RECT 79.880 109.385 81.980 109.555 ;
        RECT 79.880 109.305 80.210 109.385 ;
        RECT 80.010 108.365 80.180 109.080 ;
        RECT 80.380 109.025 81.100 109.215 ;
        RECT 81.810 109.150 81.980 109.385 ;
        RECT 81.310 108.855 81.640 109.000 ;
        RECT 80.350 108.535 81.640 108.855 ;
        RECT 81.810 108.365 81.980 108.980 ;
        RECT 80.010 108.195 81.980 108.365 ;
        RECT 82.260 108.380 82.430 109.735 ;
        RECT 82.710 109.845 84.810 110.015 ;
        RECT 82.710 109.610 82.880 109.845 ;
        RECT 84.480 109.765 84.810 109.845 ;
        RECT 83.590 109.485 84.310 109.675 ;
        RECT 82.710 108.825 82.880 109.440 ;
        RECT 83.050 109.315 83.380 109.460 ;
        RECT 83.050 108.995 84.340 109.315 ;
        RECT 84.510 108.825 84.680 109.540 ;
        RECT 82.710 108.655 84.680 108.825 ;
        RECT 84.980 108.840 86.240 110.185 ;
        RECT 86.410 109.300 87.870 110.660 ;
        RECT 88.150 110.765 90.250 110.935 ;
        RECT 88.150 110.530 88.320 110.765 ;
        RECT 89.920 110.685 90.250 110.765 ;
        RECT 89.030 110.405 89.750 110.595 ;
        RECT 88.150 109.745 88.320 110.360 ;
        RECT 88.490 110.235 88.820 110.380 ;
        RECT 88.490 109.915 89.780 110.235 ;
        RECT 89.950 109.745 90.120 110.460 ;
        RECT 88.150 109.575 90.120 109.745 ;
        RECT 86.410 109.090 88.400 109.300 ;
        RECT 86.410 109.010 87.870 109.090 ;
        RECT 77.855 108.015 79.710 108.175 ;
        RECT 77.855 107.825 80.210 108.015 ;
        RECT 73.600 106.780 74.705 107.095 ;
        RECT 75.445 106.895 77.535 107.235 ;
        RECT 71.765 106.400 72.290 106.530 ;
        RECT 72.995 106.400 73.930 106.550 ;
        RECT 71.765 106.210 73.930 106.400 ;
        RECT 71.765 106.200 72.790 106.210 ;
        RECT 71.380 105.990 72.160 106.030 ;
        RECT 70.920 105.860 72.160 105.990 ;
        RECT 70.920 105.820 71.550 105.860 ;
        RECT 70.580 105.310 71.210 105.640 ;
        RECT 69.850 104.510 70.390 105.005 ;
        RECT 70.580 104.670 70.750 105.310 ;
        RECT 71.380 105.190 71.550 105.820 ;
        RECT 71.770 105.535 72.290 105.690 ;
        RECT 72.460 105.650 72.790 106.200 ;
        RECT 74.100 106.040 74.705 106.780 ;
        RECT 73.090 105.870 74.705 106.040 ;
        RECT 71.770 105.480 72.330 105.535 ;
        RECT 72.960 105.525 73.885 105.700 ;
        RECT 72.910 105.480 73.885 105.525 ;
        RECT 71.770 105.370 73.885 105.480 ;
        RECT 74.100 105.415 74.705 105.870 ;
        RECT 76.275 106.235 77.535 106.895 ;
        RECT 79.105 107.700 80.210 107.825 ;
        RECT 79.105 106.960 79.710 107.700 ;
        RECT 80.440 107.470 80.815 108.025 ;
        RECT 81.020 107.490 81.350 108.195 ;
        RECT 82.260 108.170 82.960 108.380 ;
        RECT 82.260 107.920 82.430 108.170 ;
        RECT 83.340 107.950 83.670 108.655 ;
        RECT 81.730 107.710 82.430 107.920 ;
        RECT 83.875 107.930 84.250 108.485 ;
        RECT 84.980 108.475 86.760 108.840 ;
        RECT 84.480 108.160 86.760 108.475 ;
        RECT 79.880 107.320 80.815 107.470 ;
        RECT 81.520 107.320 82.045 107.450 ;
        RECT 79.880 107.130 82.045 107.320 ;
        RECT 81.020 107.120 82.045 107.130 ;
        RECT 82.260 107.410 82.430 107.710 ;
        RECT 82.645 107.780 83.170 107.910 ;
        RECT 83.875 107.780 84.810 107.930 ;
        RECT 82.645 107.590 84.810 107.780 ;
        RECT 82.645 107.580 83.670 107.590 ;
        RECT 82.260 107.240 83.040 107.410 ;
        RECT 79.105 106.790 80.720 106.960 ;
        RECT 79.105 106.235 79.710 106.790 ;
        RECT 79.925 106.445 80.850 106.620 ;
        RECT 81.020 106.570 81.350 107.120 ;
        RECT 82.260 106.950 82.430 107.240 ;
        RECT 81.650 106.780 82.430 106.950 ;
        RECT 81.520 106.455 82.040 106.610 ;
        RECT 79.925 106.400 80.900 106.445 ;
        RECT 81.480 106.400 82.040 106.455 ;
        RECT 79.925 106.290 82.040 106.400 ;
        RECT 76.275 106.060 76.990 106.235 ;
        RECT 79.540 106.120 79.710 106.235 ;
        RECT 80.770 106.280 82.040 106.290 ;
        RECT 82.260 106.570 82.430 106.780 ;
        RECT 82.650 106.915 83.170 107.070 ;
        RECT 83.340 107.030 83.670 107.580 ;
        RECT 84.980 107.420 86.760 108.160 ;
        RECT 83.970 107.250 86.760 107.420 ;
        RECT 84.980 107.150 86.760 107.250 ;
        RECT 86.930 108.330 87.870 109.010 ;
        RECT 88.780 108.870 89.110 109.575 ;
        RECT 89.315 108.850 89.690 109.405 ;
        RECT 90.420 109.395 90.590 111.105 ;
        RECT 92.160 110.935 92.460 111.395 ;
        RECT 92.640 111.115 93.855 111.485 ;
        RECT 90.760 110.765 92.860 110.935 ;
        RECT 90.760 110.685 91.090 110.765 ;
        RECT 90.890 109.745 91.060 110.460 ;
        RECT 91.260 110.405 91.980 110.595 ;
        RECT 92.690 110.530 92.860 110.765 ;
        RECT 93.140 110.835 93.855 111.115 ;
        RECT 95.425 112.035 96.030 112.425 ;
        RECT 96.200 112.375 97.170 112.480 ;
        RECT 97.905 112.375 98.250 112.480 ;
        RECT 96.200 112.205 98.250 112.375 ;
        RECT 98.580 112.035 98.750 112.670 ;
        RECT 101.300 112.660 101.970 112.720 ;
        RECT 102.140 112.895 102.310 113.160 ;
        RECT 102.480 113.065 103.130 113.415 ;
        RECT 103.300 113.160 103.760 113.330 ;
        RECT 103.300 112.895 103.470 113.160 ;
        RECT 104.020 113.120 104.570 113.450 ;
        RECT 104.740 113.355 104.910 113.620 ;
        RECT 105.080 113.525 105.730 113.875 ;
        RECT 105.900 113.620 106.570 113.790 ;
        RECT 105.900 113.355 106.070 113.620 ;
        RECT 106.740 113.590 108.520 114.490 ;
        RECT 108.690 114.595 110.175 114.970 ;
        RECT 108.690 114.255 111.005 114.595 ;
        RECT 108.690 113.590 110.175 114.255 ;
        RECT 106.740 113.450 106.910 113.590 ;
        RECT 104.740 113.125 106.070 113.355 ;
        RECT 106.240 113.120 106.910 113.450 ;
        RECT 107.080 113.160 107.750 113.330 ;
        RECT 104.020 112.990 104.190 113.120 ;
        RECT 102.140 112.665 103.470 112.895 ;
        RECT 103.640 112.660 104.190 112.990 ;
        RECT 106.740 112.990 106.910 113.120 ;
        RECT 104.450 112.765 106.570 112.950 ;
        RECT 99.340 112.550 100.705 112.605 ;
        RECT 99.030 112.435 101.130 112.550 ;
        RECT 99.030 112.380 99.470 112.435 ;
        RECT 99.030 112.215 99.200 112.380 ;
        RECT 100.575 112.300 101.130 112.435 ;
        RECT 95.425 111.865 97.210 112.035 ;
        RECT 97.665 111.865 98.750 112.035 ;
        RECT 95.425 111.140 96.030 111.865 ;
        RECT 96.200 111.400 98.410 111.580 ;
        RECT 96.200 111.310 97.105 111.400 ;
        RECT 97.905 111.320 98.410 111.400 ;
        RECT 95.425 110.835 96.790 111.140 ;
        RECT 97.275 111.125 97.605 111.230 ;
        RECT 98.580 111.140 98.750 111.865 ;
        RECT 99.030 111.515 99.200 112.020 ;
        RECT 99.400 111.855 99.620 112.210 ;
        RECT 99.790 112.025 100.385 112.265 ;
        RECT 99.400 111.685 100.685 111.855 ;
        RECT 99.030 111.345 100.150 111.515 ;
        RECT 93.140 110.660 93.310 110.835 ;
        RECT 95.860 110.810 96.790 110.835 ;
        RECT 96.960 110.955 98.030 111.125 ;
        RECT 95.860 110.660 96.030 110.810 ;
        RECT 92.190 110.235 92.520 110.380 ;
        RECT 91.230 109.915 92.520 110.235 ;
        RECT 92.690 109.745 92.860 110.360 ;
        RECT 90.890 109.575 92.860 109.745 ;
        RECT 89.920 109.080 91.090 109.395 ;
        RECT 88.085 108.700 88.610 108.830 ;
        RECT 89.315 108.700 90.250 108.850 ;
        RECT 88.085 108.510 90.250 108.700 ;
        RECT 88.085 108.500 89.110 108.510 ;
        RECT 86.930 108.160 88.480 108.330 ;
        RECT 86.930 107.490 87.870 108.160 ;
        RECT 88.090 107.835 88.610 107.990 ;
        RECT 88.780 107.950 89.110 108.500 ;
        RECT 90.420 108.340 90.590 109.080 ;
        RECT 91.320 108.850 91.695 109.405 ;
        RECT 91.900 108.870 92.230 109.575 ;
        RECT 93.140 109.300 93.855 110.660 ;
        RECT 92.610 109.090 93.855 109.300 ;
        RECT 93.140 109.075 93.855 109.090 ;
        RECT 95.425 110.200 96.030 110.660 ;
        RECT 96.960 110.630 97.130 110.955 ;
        RECT 96.200 110.450 97.130 110.630 ;
        RECT 97.310 110.390 97.680 110.730 ;
        RECT 97.860 110.630 98.030 110.955 ;
        RECT 98.200 111.025 98.750 111.140 ;
        RECT 99.980 111.155 100.150 111.345 ;
        RECT 100.320 111.325 100.685 111.685 ;
        RECT 100.855 111.155 101.025 112.090 ;
        RECT 98.200 110.810 99.250 111.025 ;
        RECT 98.580 110.655 99.250 110.810 ;
        RECT 99.430 110.935 99.760 111.135 ;
        RECT 99.980 110.985 101.025 111.155 ;
        RECT 101.300 112.065 101.470 112.660 ;
        RECT 104.020 112.510 104.190 112.660 ;
        RECT 106.740 112.660 107.410 112.990 ;
        RECT 107.580 112.895 107.750 113.160 ;
        RECT 107.920 113.065 108.570 113.415 ;
        RECT 108.740 113.160 109.200 113.330 ;
        RECT 108.740 112.895 108.910 113.160 ;
        RECT 109.460 112.990 110.175 113.590 ;
        RECT 107.580 112.665 108.910 112.895 ;
        RECT 109.080 112.660 110.175 112.990 ;
        RECT 111.745 112.775 112.350 116.180 ;
        RECT 101.640 112.305 103.760 112.490 ;
        RECT 104.020 112.260 104.650 112.510 ;
        RECT 104.820 112.315 105.770 112.595 ;
        RECT 106.740 112.525 106.910 112.660 ;
        RECT 106.280 112.260 106.910 112.525 ;
        RECT 107.080 112.305 109.200 112.490 ;
        RECT 101.300 111.800 101.930 112.065 ;
        RECT 102.440 111.855 103.390 112.135 ;
        RECT 104.020 112.050 104.190 112.260 ;
        RECT 104.780 112.090 106.145 112.145 ;
        RECT 103.560 111.800 104.190 112.050 ;
        RECT 97.860 110.460 98.410 110.630 ;
        RECT 98.580 110.200 98.750 110.655 ;
        RECT 99.430 110.475 99.730 110.935 ;
        RECT 99.980 110.815 100.240 110.985 ;
        RECT 101.300 110.815 101.470 111.800 ;
        RECT 102.065 111.630 103.430 111.685 ;
        RECT 101.640 111.515 103.740 111.630 ;
        RECT 101.640 111.380 102.195 111.515 ;
        RECT 103.300 111.460 103.740 111.515 ;
        RECT 99.910 110.645 100.240 110.815 ;
        RECT 100.500 110.645 101.470 110.815 ;
        RECT 90.760 108.700 91.695 108.850 ;
        RECT 92.400 108.700 92.925 108.830 ;
        RECT 90.760 108.510 92.925 108.700 ;
        RECT 91.900 108.500 92.925 108.510 ;
        RECT 93.140 108.735 94.685 109.075 ;
        RECT 89.410 108.170 91.600 108.340 ;
        RECT 88.090 107.780 88.650 107.835 ;
        RECT 89.280 107.825 90.205 108.000 ;
        RECT 89.230 107.780 90.205 107.825 ;
        RECT 88.090 107.670 90.205 107.780 ;
        RECT 88.090 107.660 89.360 107.670 ;
        RECT 88.525 107.610 89.360 107.660 ;
        RECT 90.420 107.500 90.590 108.170 ;
        RECT 90.805 107.825 91.730 108.000 ;
        RECT 91.900 107.950 92.230 108.500 ;
        RECT 93.140 108.330 93.855 108.735 ;
        RECT 92.530 108.160 93.855 108.330 ;
        RECT 92.400 107.835 92.920 107.990 ;
        RECT 90.805 107.780 91.780 107.825 ;
        RECT 92.360 107.780 92.920 107.835 ;
        RECT 90.805 107.670 92.920 107.780 ;
        RECT 91.650 107.660 92.920 107.670 ;
        RECT 91.650 107.610 92.485 107.660 ;
        RECT 86.930 107.320 88.385 107.490 ;
        RECT 89.505 107.330 91.505 107.500 ;
        RECT 93.140 107.490 93.855 108.160 ;
        RECT 86.930 107.150 87.870 107.320 ;
        RECT 82.650 106.860 83.210 106.915 ;
        RECT 83.840 106.905 84.765 107.080 ;
        RECT 83.790 106.860 84.765 106.905 ;
        RECT 82.650 106.750 84.765 106.860 ;
        RECT 82.650 106.740 83.920 106.750 ;
        RECT 83.085 106.690 83.920 106.740 ;
        RECT 84.980 106.580 85.150 107.150 ;
        RECT 82.260 106.400 82.945 106.570 ;
        RECT 84.065 106.410 85.150 106.580 ;
        RECT 87.700 106.980 87.870 107.150 ;
        RECT 90.420 106.980 90.590 107.330 ;
        RECT 92.625 107.320 93.855 107.490 ;
        RECT 93.140 106.980 93.855 107.320 ;
        RECT 95.425 107.255 96.465 110.200 ;
        RECT 98.035 108.840 98.750 110.200 ;
        RECT 99.030 110.305 101.130 110.475 ;
        RECT 99.030 110.070 99.200 110.305 ;
        RECT 100.800 110.225 101.130 110.305 ;
        RECT 99.910 109.945 100.630 110.135 ;
        RECT 99.030 109.285 99.200 109.900 ;
        RECT 99.370 109.775 99.700 109.920 ;
        RECT 99.370 109.455 100.660 109.775 ;
        RECT 100.830 109.285 101.000 110.000 ;
        RECT 99.030 109.115 101.000 109.285 ;
        RECT 101.300 109.895 101.470 110.645 ;
        RECT 101.745 110.235 101.915 111.170 ;
        RECT 102.385 111.105 102.980 111.345 ;
        RECT 103.570 111.295 103.740 111.460 ;
        RECT 103.150 110.935 103.370 111.290 ;
        RECT 102.085 110.765 103.370 110.935 ;
        RECT 102.085 110.405 102.450 110.765 ;
        RECT 103.570 110.595 103.740 111.100 ;
        RECT 102.620 110.425 103.740 110.595 ;
        RECT 104.020 110.565 104.190 111.800 ;
        RECT 104.470 111.975 106.570 112.090 ;
        RECT 104.470 111.920 104.910 111.975 ;
        RECT 104.470 111.755 104.640 111.920 ;
        RECT 106.015 111.840 106.570 111.975 ;
        RECT 106.740 112.065 106.910 112.260 ;
        RECT 104.470 111.055 104.640 111.560 ;
        RECT 104.840 111.395 105.060 111.750 ;
        RECT 105.230 111.565 105.825 111.805 ;
        RECT 106.740 111.800 107.370 112.065 ;
        RECT 107.880 111.855 108.830 112.135 ;
        RECT 109.460 112.050 110.175 112.660 ;
        RECT 110.495 112.425 112.350 112.775 ;
        RECT 109.000 111.800 110.175 112.050 ;
        RECT 104.840 111.225 106.125 111.395 ;
        RECT 104.470 110.885 105.590 111.055 ;
        RECT 105.420 110.695 105.590 110.885 ;
        RECT 105.760 110.865 106.125 111.225 ;
        RECT 106.295 110.695 106.465 111.630 ;
        RECT 102.620 110.235 102.790 110.425 ;
        RECT 101.745 110.065 102.790 110.235 ;
        RECT 102.530 109.895 102.790 110.065 ;
        RECT 103.010 110.015 103.340 110.215 ;
        RECT 104.020 110.195 104.690 110.565 ;
        RECT 104.870 110.475 105.200 110.675 ;
        RECT 105.420 110.525 106.465 110.695 ;
        RECT 104.020 110.105 104.190 110.195 ;
        RECT 101.300 109.725 102.270 109.895 ;
        RECT 102.530 109.725 102.860 109.895 ;
        RECT 98.035 108.630 99.280 108.840 ;
        RECT 98.035 108.615 98.750 108.630 ;
        RECT 97.205 108.275 98.750 108.615 ;
        RECT 99.660 108.410 99.990 109.115 ;
        RECT 100.195 108.390 100.570 108.945 ;
        RECT 101.300 108.935 101.470 109.725 ;
        RECT 103.040 109.555 103.340 110.015 ;
        RECT 103.520 109.735 104.190 110.105 ;
        RECT 104.870 110.015 105.170 110.475 ;
        RECT 105.420 110.355 105.680 110.525 ;
        RECT 106.740 110.355 106.910 111.800 ;
        RECT 107.505 111.630 108.870 111.685 ;
        RECT 107.080 111.515 109.180 111.630 ;
        RECT 107.080 111.380 107.635 111.515 ;
        RECT 108.740 111.460 109.180 111.515 ;
        RECT 105.350 110.185 105.680 110.355 ;
        RECT 105.940 110.185 106.910 110.355 ;
        RECT 101.640 109.385 103.740 109.555 ;
        RECT 101.640 109.305 101.970 109.385 ;
        RECT 100.800 108.620 101.470 108.935 ;
        RECT 80.770 106.230 81.605 106.280 ;
        RECT 79.540 106.060 80.625 106.120 ;
        RECT 82.260 106.110 82.430 106.400 ;
        RECT 76.275 105.540 78.280 106.060 ;
        RECT 78.450 105.950 80.625 106.060 ;
        RECT 81.745 106.060 82.430 106.110 ;
        RECT 84.980 106.060 85.150 106.410 ;
        RECT 71.770 105.360 73.040 105.370 ;
        RECT 72.205 105.310 73.040 105.360 ;
        RECT 74.100 105.200 75.955 105.415 ;
        RECT 71.380 105.080 72.065 105.190 ;
        RECT 70.920 105.020 72.065 105.080 ;
        RECT 73.185 105.065 75.955 105.200 ;
        RECT 73.185 105.030 74.705 105.065 ;
        RECT 70.920 104.910 71.550 105.020 ;
        RECT 71.380 104.680 71.550 104.910 ;
        RECT 74.100 104.680 74.705 105.030 ;
        RECT 69.850 104.450 70.020 104.510 ;
        RECT 70.580 104.340 71.210 104.670 ;
        RECT 69.000 104.170 69.680 104.195 ;
        RECT 69.000 103.960 70.870 104.170 ;
        RECT 71.040 103.790 71.210 104.340 ;
        RECT 68.660 103.480 69.895 103.790 ;
        RECT 64.360 102.990 65.030 103.160 ;
        RECT 65.200 103.065 65.640 103.235 ;
        RECT 62.785 102.645 64.190 102.815 ;
        RECT 60.500 102.295 62.045 102.635 ;
        RECT 60.500 98.875 61.215 102.295 ;
        RECT 62.785 100.815 63.390 102.645 ;
        RECT 64.360 102.240 64.530 102.990 ;
        RECT 65.940 102.960 66.610 103.295 ;
        RECT 65.940 102.895 66.110 102.960 ;
        RECT 66.780 102.945 67.350 103.300 ;
        RECT 67.520 102.975 67.980 103.300 ;
        RECT 64.700 102.410 65.260 102.820 ;
        RECT 65.430 102.580 66.110 102.895 ;
        RECT 67.470 102.775 67.640 102.780 ;
        RECT 66.330 102.590 66.850 102.760 ;
        RECT 65.940 102.390 66.110 102.580 ;
        RECT 65.430 102.240 65.770 102.350 ;
        RECT 64.360 102.060 65.770 102.240 ;
        RECT 65.940 102.060 66.510 102.390 ;
        RECT 64.185 101.700 64.530 102.060 ;
        RECT 65.940 101.890 66.110 102.060 ;
        RECT 66.680 101.890 66.850 102.590 ;
        RECT 67.020 102.065 67.640 102.775 ;
        RECT 64.700 101.695 65.260 101.890 ;
        RECT 65.090 101.690 65.260 101.695 ;
        RECT 65.430 101.650 66.110 101.890 ;
        RECT 66.330 101.720 66.850 101.890 ;
        RECT 65.940 101.550 66.110 101.650 ;
        RECT 61.535 100.465 63.390 100.815 ;
        RECT 62.785 99.480 63.390 100.465 ;
        RECT 63.560 101.010 64.230 101.260 ;
        RECT 64.400 101.050 65.300 101.460 ;
        RECT 65.940 101.220 66.510 101.550 ;
        RECT 65.470 101.170 66.510 101.220 ;
        RECT 66.680 101.320 66.850 101.720 ;
        RECT 67.020 101.490 67.350 101.895 ;
        RECT 67.810 101.875 67.980 102.975 ;
        RECT 67.520 101.705 67.980 101.875 ;
        RECT 67.520 101.320 67.690 101.705 ;
        RECT 68.150 101.640 68.440 103.300 ;
        RECT 68.660 102.770 68.830 103.480 ;
        RECT 70.065 103.475 70.700 103.790 ;
        RECT 70.870 103.480 71.210 103.790 ;
        RECT 71.380 104.390 72.275 104.680 ;
        RECT 72.935 104.390 74.705 104.680 ;
        RECT 71.380 104.220 71.550 104.390 ;
        RECT 74.100 104.220 74.705 104.390 ;
        RECT 71.380 103.470 72.840 104.220 ;
        RECT 73.010 103.475 74.705 104.220 ;
        RECT 76.275 104.850 77.740 105.540 ;
        RECT 78.450 105.370 79.710 105.950 ;
        RECT 81.745 105.940 83.720 106.060 ;
        RECT 77.910 104.850 79.710 105.370 ;
        RECT 76.275 104.680 76.990 104.850 ;
        RECT 79.540 104.680 79.710 104.850 ;
        RECT 82.260 105.540 83.720 105.940 ;
        RECT 82.260 104.850 83.180 105.540 ;
        RECT 83.890 105.370 85.150 106.060 ;
        RECT 83.350 104.850 85.150 105.370 ;
        RECT 85.370 104.860 85.660 106.520 ;
        RECT 85.830 106.195 86.290 106.520 ;
        RECT 85.830 105.095 86.000 106.195 ;
        RECT 86.460 106.165 87.030 106.520 ;
        RECT 87.700 106.515 89.160 106.980 ;
        RECT 87.200 106.230 89.160 106.515 ;
        RECT 87.200 106.180 88.640 106.230 ;
        RECT 86.170 105.995 86.340 106.000 ;
        RECT 86.170 105.285 86.790 105.995 ;
        RECT 86.960 105.810 87.480 105.980 ;
        RECT 85.830 104.925 86.290 105.095 ;
        RECT 82.260 104.680 82.430 104.850 ;
        RECT 84.980 104.690 85.150 104.850 ;
        RECT 84.980 104.680 85.950 104.690 ;
        RECT 76.275 104.390 77.715 104.680 ;
        RECT 78.375 104.390 80.915 104.680 ;
        RECT 81.430 104.390 83.155 104.680 ;
        RECT 83.815 104.410 85.950 104.680 ;
        RECT 86.120 104.540 86.290 104.925 ;
        RECT 86.460 104.710 86.790 105.115 ;
        RECT 86.960 105.110 87.130 105.810 ;
        RECT 87.700 105.610 88.640 106.180 ;
        RECT 89.330 106.060 91.680 106.980 ;
        RECT 91.850 106.230 93.855 106.980 ;
        RECT 94.175 106.905 96.465 107.255 ;
        RECT 87.300 105.310 88.640 105.610 ;
        RECT 88.810 105.310 92.200 106.060 ;
        RECT 92.370 105.315 93.855 106.230 ;
        RECT 95.425 106.795 96.465 106.905 ;
        RECT 98.035 107.870 98.750 108.275 ;
        RECT 98.965 108.240 99.490 108.370 ;
        RECT 100.195 108.240 101.130 108.390 ;
        RECT 98.965 108.050 101.130 108.240 ;
        RECT 98.965 108.040 99.990 108.050 ;
        RECT 98.035 107.700 99.360 107.870 ;
        RECT 98.035 107.030 98.750 107.700 ;
        RECT 98.970 107.375 99.490 107.530 ;
        RECT 99.660 107.490 99.990 108.040 ;
        RECT 101.300 108.015 101.470 108.620 ;
        RECT 101.770 108.365 101.940 109.080 ;
        RECT 102.140 109.025 102.860 109.215 ;
        RECT 103.570 109.150 103.740 109.385 ;
        RECT 103.070 108.855 103.400 109.000 ;
        RECT 102.110 108.535 103.400 108.855 ;
        RECT 103.570 108.365 103.740 108.980 ;
        RECT 101.770 108.195 103.740 108.365 ;
        RECT 104.020 108.380 104.190 109.735 ;
        RECT 104.470 109.845 106.570 110.015 ;
        RECT 104.470 109.610 104.640 109.845 ;
        RECT 106.240 109.765 106.570 109.845 ;
        RECT 106.740 109.895 106.910 110.185 ;
        RECT 107.185 110.235 107.355 111.170 ;
        RECT 107.825 111.105 108.420 111.345 ;
        RECT 109.010 111.295 109.180 111.460 ;
        RECT 108.590 110.935 108.810 111.290 ;
        RECT 107.525 110.765 108.810 110.935 ;
        RECT 107.525 110.405 107.890 110.765 ;
        RECT 109.010 110.595 109.180 111.100 ;
        RECT 108.060 110.425 109.180 110.595 ;
        RECT 109.460 110.835 110.175 111.800 ;
        RECT 111.745 110.835 112.350 112.425 ;
        RECT 109.460 110.660 109.630 110.835 ;
        RECT 112.180 110.660 112.350 110.835 ;
        RECT 108.060 110.235 108.230 110.425 ;
        RECT 107.185 110.065 108.230 110.235 ;
        RECT 107.970 109.895 108.230 110.065 ;
        RECT 108.450 110.015 108.780 110.215 ;
        RECT 109.460 110.105 110.175 110.660 ;
        RECT 106.740 109.725 107.710 109.895 ;
        RECT 107.970 109.725 108.300 109.895 ;
        RECT 105.350 109.485 106.070 109.675 ;
        RECT 104.470 108.825 104.640 109.440 ;
        RECT 104.810 109.315 105.140 109.460 ;
        RECT 104.810 108.995 106.100 109.315 ;
        RECT 106.270 108.825 106.440 109.540 ;
        RECT 104.470 108.655 106.440 108.825 ;
        RECT 101.300 107.880 101.970 108.015 ;
        RECT 100.290 107.710 101.970 107.880 ;
        RECT 101.300 107.700 101.970 107.710 ;
        RECT 98.970 107.320 99.530 107.375 ;
        RECT 100.160 107.365 101.085 107.540 ;
        RECT 100.110 107.320 101.085 107.365 ;
        RECT 98.970 107.210 101.085 107.320 ;
        RECT 98.970 107.200 100.240 107.210 ;
        RECT 99.405 107.150 100.240 107.200 ;
        RECT 101.300 107.040 101.470 107.700 ;
        RECT 102.200 107.470 102.575 108.025 ;
        RECT 102.780 107.490 103.110 108.195 ;
        RECT 104.020 108.170 104.720 108.380 ;
        RECT 104.020 107.920 104.190 108.170 ;
        RECT 105.100 107.950 105.430 108.655 ;
        RECT 103.490 107.710 104.190 107.920 ;
        RECT 105.635 107.930 106.010 108.485 ;
        RECT 106.740 108.475 106.910 109.725 ;
        RECT 108.480 109.555 108.780 110.015 ;
        RECT 108.960 109.735 110.175 110.105 ;
        RECT 107.080 109.385 109.180 109.555 ;
        RECT 107.080 109.305 107.410 109.385 ;
        RECT 106.240 108.160 106.910 108.475 ;
        RECT 107.210 108.365 107.380 109.080 ;
        RECT 107.580 109.025 108.300 109.215 ;
        RECT 109.010 109.150 109.180 109.385 ;
        RECT 109.460 109.075 110.175 109.735 ;
        RECT 108.510 108.855 108.840 109.000 ;
        RECT 107.550 108.535 108.840 108.855 ;
        RECT 109.010 108.365 109.180 108.980 ;
        RECT 107.210 108.195 109.180 108.365 ;
        RECT 109.460 108.735 111.005 109.075 ;
        RECT 106.740 108.015 106.910 108.160 ;
        RECT 101.640 107.320 102.575 107.470 ;
        RECT 103.280 107.320 103.805 107.450 ;
        RECT 101.640 107.130 103.805 107.320 ;
        RECT 98.035 106.860 99.265 107.030 ;
        RECT 100.385 106.960 101.470 107.040 ;
        RECT 102.780 107.120 103.805 107.130 ;
        RECT 104.020 107.410 104.190 107.710 ;
        RECT 104.405 107.780 104.930 107.910 ;
        RECT 105.635 107.780 106.570 107.930 ;
        RECT 104.405 107.590 106.570 107.780 ;
        RECT 106.740 107.700 107.410 108.015 ;
        RECT 104.405 107.580 105.430 107.590 ;
        RECT 104.020 107.240 104.800 107.410 ;
        RECT 100.385 106.870 102.480 106.960 ;
        RECT 95.425 106.445 97.715 106.795 ;
        RECT 98.035 106.520 98.750 106.860 ;
        RECT 101.300 106.790 102.480 106.870 ;
        RECT 101.300 106.520 101.470 106.790 ;
        RECT 95.425 105.315 96.465 106.445 ;
        RECT 92.370 105.310 93.310 105.315 ;
        RECT 87.300 105.280 87.870 105.310 ;
        RECT 86.960 104.940 87.480 105.110 ;
        RECT 86.960 104.540 87.130 104.940 ;
        RECT 87.700 104.770 87.870 105.280 ;
        RECT 83.815 104.390 85.150 104.410 ;
        RECT 76.275 104.220 76.990 104.390 ;
        RECT 79.540 104.220 79.710 104.390 ;
        RECT 76.275 103.475 77.535 104.220 ;
        RECT 71.380 103.270 72.320 103.470 ;
        RECT 73.010 103.300 74.270 103.475 ;
        RECT 76.820 103.300 77.535 103.475 ;
        RECT 69.000 102.940 69.620 103.270 ;
        RECT 69.850 102.975 70.470 103.265 ;
        RECT 70.640 102.940 72.320 103.270 ;
        RECT 68.660 102.600 69.280 102.770 ;
        RECT 68.660 101.470 68.830 102.600 ;
        RECT 69.450 102.430 69.620 102.940 ;
        RECT 69.000 102.100 69.620 102.430 ;
        RECT 69.850 102.390 70.470 102.805 ;
        RECT 71.380 102.550 72.320 102.940 ;
        RECT 72.490 102.550 74.705 103.300 ;
        RECT 70.640 102.220 70.830 102.445 ;
        RECT 69.790 102.050 70.830 102.220 ;
        RECT 69.790 101.930 69.960 102.050 ;
        RECT 71.380 102.010 71.550 102.550 ;
        RECT 69.000 101.760 69.960 101.930 ;
        RECT 69.000 101.680 69.570 101.760 ;
        RECT 65.470 101.050 66.110 101.170 ;
        RECT 66.680 101.150 67.690 101.320 ;
        RECT 67.860 101.190 68.830 101.470 ;
        RECT 63.560 100.420 63.730 101.010 ;
        RECT 64.400 100.840 64.610 101.050 ;
        RECT 65.120 100.880 65.300 101.050 ;
        RECT 63.900 100.590 64.610 100.840 ;
        RECT 63.560 99.650 64.240 100.420 ;
        RECT 64.780 100.350 64.950 100.840 ;
        RECT 62.785 99.175 63.890 99.480 ;
        RECT 62.785 98.875 63.390 99.175 ;
        RECT 64.070 99.005 64.240 99.650 ;
        RECT 60.500 97.270 60.670 98.875 ;
        RECT 63.220 98.585 63.390 98.875 ;
        RECT 63.560 98.755 64.240 99.005 ;
        RECT 63.220 98.335 63.890 98.585 ;
        RECT 63.220 97.780 63.390 98.335 ;
        RECT 64.070 98.165 64.240 98.755 ;
        RECT 63.560 97.955 64.240 98.165 ;
        RECT 64.410 100.180 64.950 100.350 ;
        RECT 65.120 100.550 65.380 100.880 ;
        RECT 63.560 97.850 63.900 97.955 ;
        RECT 64.410 97.785 64.580 100.180 ;
        RECT 65.120 100.020 65.300 100.550 ;
        RECT 65.940 100.535 66.110 101.050 ;
        RECT 67.020 101.045 67.350 101.150 ;
        RECT 68.660 101.075 68.830 101.190 ;
        RECT 66.440 100.875 66.785 100.980 ;
        RECT 67.520 100.875 68.490 100.980 ;
        RECT 66.440 100.705 68.490 100.875 ;
        RECT 68.660 100.745 69.190 101.075 ;
        RECT 69.360 100.990 69.570 101.680 ;
        RECT 70.140 101.570 70.470 101.880 ;
        RECT 71.000 101.815 71.550 102.010 ;
        RECT 71.000 101.680 72.020 101.815 ;
        RECT 71.380 101.645 72.020 101.680 ;
        RECT 72.190 101.715 73.420 101.885 ;
        RECT 73.600 101.860 73.930 101.885 ;
        RECT 69.740 101.400 70.810 101.570 ;
        RECT 69.740 101.160 69.910 101.400 ;
        RECT 70.140 101.035 70.470 101.230 ;
        RECT 70.640 101.160 70.810 101.400 ;
        RECT 69.360 100.820 69.970 100.990 ;
        RECT 68.660 100.535 68.830 100.745 ;
        RECT 69.800 100.605 69.970 100.820 ;
        RECT 70.140 100.775 70.430 101.035 ;
        RECT 71.380 100.975 71.550 101.645 ;
        RECT 72.190 101.475 72.370 101.715 ;
        RECT 71.720 101.145 72.370 101.475 ;
        RECT 71.380 100.925 72.020 100.975 ;
        RECT 70.600 100.805 72.020 100.925 ;
        RECT 70.600 100.725 71.550 100.805 ;
        RECT 65.940 100.380 67.025 100.535 ;
        RECT 65.470 100.365 67.025 100.380 ;
        RECT 67.480 100.365 68.830 100.535 ;
        RECT 65.470 100.210 66.110 100.365 ;
        RECT 65.090 99.850 65.300 100.020 ;
        RECT 64.750 98.985 64.950 99.655 ;
        RECT 65.120 99.520 65.300 99.850 ;
        RECT 65.120 99.190 65.380 99.520 ;
        RECT 65.550 98.965 65.770 99.945 ;
        RECT 60.840 97.440 61.470 97.780 ;
        RECT 60.500 97.100 61.130 97.270 ;
        RECT 60.500 95.480 60.670 97.100 ;
        RECT 61.300 96.930 61.470 97.440 ;
        RECT 61.660 97.020 61.910 97.780 ;
        RECT 62.080 97.520 63.390 97.780 ;
        RECT 62.080 97.020 63.050 97.350 ;
        RECT 60.840 96.680 61.470 96.930 ;
        RECT 60.840 96.090 61.050 96.680 ;
        RECT 60.840 95.760 61.070 96.090 ;
        RECT 61.240 95.930 61.490 96.510 ;
        RECT 61.660 96.100 61.910 96.850 ;
        RECT 62.080 96.510 62.250 97.020 ;
        RECT 63.220 96.850 63.390 97.520 ;
        RECT 62.420 96.680 63.390 96.850 ;
        RECT 62.080 96.180 63.050 96.510 ;
        RECT 63.220 96.385 63.390 96.680 ;
        RECT 63.560 97.395 63.890 97.645 ;
        RECT 64.070 97.615 64.580 97.785 ;
        RECT 63.560 96.805 63.730 97.395 ;
        RECT 64.070 97.225 64.240 97.615 ;
        RECT 64.750 97.445 64.950 98.795 ;
        RECT 65.120 98.715 65.770 98.965 ;
        RECT 65.940 98.880 66.110 100.210 ;
        RECT 68.660 100.130 68.830 100.365 ;
        RECT 69.040 100.300 69.630 100.555 ;
        RECT 68.660 99.795 69.210 100.130 ;
        RECT 69.460 100.085 69.630 100.300 ;
        RECT 69.800 100.275 70.390 100.605 ;
        RECT 70.580 100.225 71.150 100.555 ;
        RECT 70.580 100.085 70.750 100.225 ;
        RECT 69.460 99.855 70.750 100.085 ;
        RECT 71.380 100.135 71.550 100.725 ;
        RECT 72.190 100.635 72.370 101.145 ;
        RECT 72.540 101.300 72.740 101.460 ;
        RECT 72.540 101.130 73.080 101.300 ;
        RECT 71.720 100.305 72.370 100.635 ;
        RECT 72.540 100.465 72.740 100.960 ;
        RECT 72.910 100.295 73.080 101.130 ;
        RECT 71.380 100.050 72.020 100.135 ;
        RECT 70.920 99.965 72.020 100.050 ;
        RECT 72.540 100.125 73.080 100.295 ;
        RECT 73.250 100.595 73.420 101.715 ;
        RECT 73.590 101.690 73.930 101.860 ;
        RECT 73.600 101.605 73.930 101.690 ;
        RECT 74.100 101.435 74.705 102.550 ;
        RECT 76.275 102.635 77.535 103.300 ;
        RECT 79.105 103.735 79.710 104.220 ;
        RECT 79.880 104.050 81.930 104.220 ;
        RECT 79.880 103.945 80.850 104.050 ;
        RECT 81.585 103.945 81.930 104.050 ;
        RECT 81.020 103.775 81.350 103.880 ;
        RECT 79.105 103.455 80.510 103.735 ;
        RECT 80.680 103.605 81.690 103.775 ;
        RECT 82.260 103.755 82.430 104.390 ;
        RECT 76.275 102.295 78.365 102.635 ;
        RECT 76.275 101.715 77.535 102.295 ;
        RECT 73.600 101.185 74.705 101.435 ;
        RECT 75.445 101.375 77.535 101.715 ;
        RECT 73.600 100.940 73.930 101.015 ;
        RECT 73.590 100.770 73.930 100.940 ;
        RECT 73.600 100.765 73.930 100.770 ;
        RECT 73.250 100.345 73.590 100.595 ;
        RECT 70.190 99.850 70.360 99.855 ;
        RECT 70.920 99.795 71.550 99.965 ;
        RECT 68.660 99.620 68.830 99.795 ;
        RECT 71.380 99.620 71.550 99.795 ;
        RECT 66.920 99.345 68.310 99.620 ;
        RECT 66.315 99.280 68.310 99.345 ;
        RECT 66.315 99.100 67.090 99.280 ;
        RECT 65.120 98.205 65.300 98.715 ;
        RECT 65.940 98.545 66.645 98.880 ;
        RECT 65.470 98.375 66.645 98.545 ;
        RECT 66.920 98.390 67.090 99.100 ;
        RECT 67.465 98.530 67.655 99.110 ;
        RECT 67.900 99.105 68.310 99.280 ;
        RECT 68.660 98.930 69.920 99.620 ;
        RECT 70.090 99.195 71.550 99.620 ;
        RECT 71.720 99.365 72.370 99.695 ;
        RECT 70.090 99.100 72.020 99.195 ;
        RECT 70.630 99.025 72.020 99.100 ;
        RECT 68.660 98.870 70.460 98.930 ;
        RECT 67.900 98.700 70.460 98.870 ;
        RECT 65.940 98.370 66.645 98.375 ;
        RECT 65.120 97.875 65.770 98.205 ;
        RECT 65.940 97.605 66.110 98.370 ;
        RECT 67.465 98.360 68.490 98.530 ;
        RECT 66.280 98.000 67.810 98.190 ;
        RECT 63.900 96.975 64.240 97.225 ;
        RECT 63.560 96.800 63.890 96.805 ;
        RECT 63.560 96.630 63.900 96.800 ;
        RECT 63.560 96.555 63.890 96.630 ;
        RECT 62.080 95.930 62.250 96.180 ;
        RECT 63.220 96.135 63.890 96.385 ;
        RECT 63.220 96.010 63.390 96.135 ;
        RECT 61.240 95.650 62.250 95.930 ;
        RECT 62.420 95.755 63.390 96.010 ;
        RECT 63.220 95.480 63.390 95.755 ;
        RECT 63.560 95.880 63.890 95.965 ;
        RECT 63.560 95.710 63.900 95.880 ;
        RECT 64.070 95.855 64.240 96.975 ;
        RECT 64.410 97.275 64.950 97.445 ;
        RECT 65.470 97.435 66.110 97.605 ;
        RECT 66.280 97.555 67.440 97.830 ;
        RECT 66.450 97.550 66.620 97.555 ;
        RECT 64.410 96.440 64.580 97.275 ;
        RECT 64.750 96.610 64.950 97.105 ;
        RECT 65.120 96.935 65.770 97.265 ;
        RECT 64.410 96.270 64.950 96.440 ;
        RECT 64.750 96.110 64.950 96.270 ;
        RECT 65.120 96.425 65.300 96.935 ;
        RECT 65.940 96.765 66.110 97.435 ;
        RECT 66.280 97.010 66.645 97.365 ;
        RECT 67.640 97.350 67.810 98.000 ;
        RECT 66.840 97.180 67.810 97.350 ;
        RECT 67.980 97.010 68.150 97.965 ;
        RECT 66.280 96.840 68.150 97.010 ;
        RECT 66.280 96.835 66.850 96.840 ;
        RECT 65.470 96.595 66.110 96.765 ;
        RECT 65.120 96.095 65.770 96.425 ;
        RECT 65.940 96.410 66.110 96.595 ;
        RECT 65.120 95.855 65.300 96.095 ;
        RECT 65.940 96.080 66.510 96.410 ;
        RECT 66.680 96.250 66.850 96.835 ;
        RECT 68.320 96.670 68.490 98.360 ;
        RECT 67.020 96.500 68.490 96.670 ;
        RECT 68.660 98.410 70.460 98.700 ;
        RECT 70.630 98.410 71.550 99.025 ;
        RECT 72.190 98.855 72.370 99.365 ;
        RECT 68.660 97.785 68.830 98.410 ;
        RECT 71.380 98.225 71.550 98.410 ;
        RECT 69.000 97.955 69.610 98.215 ;
        RECT 68.660 97.455 69.190 97.785 ;
        RECT 68.660 96.850 68.830 97.455 ;
        RECT 69.360 97.275 69.610 97.955 ;
        RECT 69.000 97.105 69.610 97.275 ;
        RECT 68.660 96.680 69.270 96.850 ;
        RECT 67.020 96.475 67.350 96.500 ;
        RECT 68.660 96.330 68.830 96.680 ;
        RECT 69.440 96.510 69.610 97.105 ;
        RECT 66.680 96.080 67.350 96.250 ;
        RECT 67.520 96.160 68.830 96.330 ;
        RECT 65.940 95.925 66.110 96.080 ;
        RECT 67.020 95.995 67.350 96.080 ;
        RECT 63.560 95.685 63.890 95.710 ;
        RECT 64.070 95.685 65.300 95.855 ;
        RECT 65.470 95.755 66.110 95.925 ;
        RECT 65.940 95.480 66.110 95.755 ;
        RECT 66.280 95.825 66.850 95.910 ;
        RECT 67.520 95.825 68.490 95.990 ;
        RECT 66.280 95.655 68.490 95.825 ;
        RECT 60.500 93.830 61.960 95.480 ;
        RECT 62.130 94.790 64.480 95.480 ;
        RECT 64.650 95.020 66.110 95.480 ;
        RECT 68.660 95.020 68.830 96.160 ;
        RECT 69.000 96.180 69.610 96.510 ;
        RECT 69.790 97.680 70.430 98.180 ;
        RECT 70.600 97.930 71.550 98.225 ;
        RECT 69.790 96.720 69.970 97.680 ;
        RECT 70.140 96.900 70.470 97.510 ;
        RECT 70.680 97.025 71.210 97.370 ;
        RECT 71.380 97.360 71.550 97.930 ;
        RECT 71.720 98.605 72.370 98.855 ;
        RECT 72.540 98.775 72.740 100.125 ;
        RECT 73.250 99.955 73.420 100.345 ;
        RECT 73.760 100.175 73.930 100.765 ;
        RECT 72.910 99.785 73.420 99.955 ;
        RECT 73.600 99.925 73.930 100.175 ;
        RECT 74.100 99.895 74.705 101.185 ;
        RECT 71.720 97.625 71.940 98.605 ;
        RECT 72.110 98.050 72.370 98.380 ;
        RECT 71.380 97.190 72.020 97.360 ;
        RECT 69.790 96.395 70.390 96.720 ;
        RECT 70.220 96.390 70.390 96.395 ;
        RECT 69.000 95.540 69.180 96.180 ;
        RECT 70.680 96.030 70.850 97.025 ;
        RECT 71.380 96.565 71.550 97.190 ;
        RECT 72.190 97.020 72.370 98.050 ;
        RECT 72.540 97.915 72.740 98.585 ;
        RECT 72.910 97.390 73.080 99.785 ;
        RECT 73.590 99.615 73.930 99.720 ;
        RECT 72.110 96.690 72.370 97.020 ;
        RECT 72.540 97.220 73.080 97.390 ;
        RECT 73.250 99.405 73.930 99.615 ;
        RECT 74.100 99.545 75.955 99.895 ;
        RECT 73.250 98.815 73.420 99.405 ;
        RECT 74.100 99.235 74.705 99.545 ;
        RECT 73.600 98.985 74.705 99.235 ;
        RECT 73.250 98.565 73.930 98.815 ;
        RECT 73.250 97.920 73.420 98.565 ;
        RECT 74.100 98.395 74.705 98.985 ;
        RECT 73.600 98.090 74.705 98.395 ;
        RECT 74.100 97.955 74.705 98.090 ;
        RECT 76.275 98.875 77.535 101.375 ;
        RECT 79.105 101.435 79.710 103.455 ;
        RECT 79.930 102.090 80.220 103.285 ;
        RECT 80.680 103.275 80.850 103.605 ;
        RECT 80.390 103.105 80.850 103.275 ;
        RECT 80.390 102.440 80.560 103.105 ;
        RECT 81.020 102.835 81.350 103.435 ;
        RECT 80.730 102.610 81.350 102.835 ;
        RECT 81.520 103.205 81.690 103.605 ;
        RECT 81.860 103.375 82.430 103.755 ;
        RECT 81.520 103.035 82.040 103.205 ;
        RECT 80.390 102.110 80.850 102.440 ;
        RECT 81.020 102.090 81.350 102.440 ;
        RECT 81.520 102.365 81.690 103.035 ;
        RECT 82.260 102.865 82.430 103.375 ;
        RECT 84.980 103.755 85.150 104.390 ;
        RECT 86.120 104.370 87.130 104.540 ;
        RECT 87.300 104.680 87.870 104.770 ;
        RECT 90.420 104.680 90.590 105.310 ;
        RECT 87.300 104.390 88.595 104.680 ;
        RECT 89.255 104.670 90.590 104.680 ;
        RECT 93.140 104.680 93.310 105.310 ;
        RECT 95.860 104.855 96.465 105.315 ;
        RECT 98.035 105.770 100.040 106.520 ;
        RECT 100.210 106.120 101.470 106.520 ;
        RECT 101.685 106.445 102.610 106.620 ;
        RECT 102.780 106.570 103.110 107.120 ;
        RECT 104.020 106.950 104.190 107.240 ;
        RECT 103.410 106.780 104.190 106.950 ;
        RECT 103.280 106.455 103.800 106.610 ;
        RECT 101.685 106.400 102.660 106.445 ;
        RECT 103.240 106.400 103.800 106.455 ;
        RECT 101.685 106.290 103.800 106.400 ;
        RECT 102.530 106.280 103.800 106.290 ;
        RECT 104.020 106.570 104.190 106.780 ;
        RECT 104.410 106.915 104.930 107.070 ;
        RECT 105.100 107.030 105.430 107.580 ;
        RECT 106.740 107.420 106.910 107.700 ;
        RECT 107.640 107.470 108.015 108.025 ;
        RECT 108.220 107.490 108.550 108.195 ;
        RECT 109.460 107.920 110.175 108.735 ;
        RECT 108.930 107.710 110.175 107.920 ;
        RECT 105.730 107.250 106.910 107.420 ;
        RECT 104.410 106.860 104.970 106.915 ;
        RECT 105.600 106.905 106.525 107.080 ;
        RECT 105.550 106.860 106.525 106.905 ;
        RECT 104.410 106.750 106.525 106.860 ;
        RECT 106.740 106.960 106.910 107.250 ;
        RECT 107.080 107.320 108.015 107.470 ;
        RECT 108.720 107.320 109.245 107.450 ;
        RECT 107.080 107.130 109.245 107.320 ;
        RECT 108.220 107.120 109.245 107.130 ;
        RECT 106.740 106.790 107.920 106.960 ;
        RECT 104.410 106.740 105.680 106.750 ;
        RECT 104.845 106.690 105.680 106.740 ;
        RECT 106.740 106.580 106.910 106.790 ;
        RECT 104.020 106.400 104.705 106.570 ;
        RECT 105.825 106.410 106.910 106.580 ;
        RECT 102.530 106.230 103.365 106.280 ;
        RECT 100.210 105.950 102.385 106.120 ;
        RECT 104.020 106.110 104.190 106.400 ;
        RECT 103.505 106.060 104.190 106.110 ;
        RECT 106.740 106.120 106.910 106.410 ;
        RECT 107.125 106.445 108.050 106.620 ;
        RECT 108.220 106.570 108.550 107.120 ;
        RECT 109.460 106.950 110.175 107.710 ;
        RECT 111.745 107.255 112.350 110.660 ;
        RECT 108.850 106.780 110.175 106.950 ;
        RECT 110.495 106.905 112.350 107.255 ;
        RECT 108.720 106.455 109.240 106.610 ;
        RECT 107.125 106.400 108.100 106.445 ;
        RECT 108.680 106.400 109.240 106.455 ;
        RECT 107.125 106.290 109.240 106.400 ;
        RECT 107.970 106.280 109.240 106.290 ;
        RECT 107.970 106.230 108.805 106.280 ;
        RECT 106.740 106.060 107.825 106.120 ;
        RECT 109.460 106.110 110.175 106.780 ;
        RECT 98.035 104.855 99.520 105.770 ;
        RECT 100.210 105.600 101.470 105.950 ;
        RECT 103.505 105.940 105.480 106.060 ;
        RECT 95.860 104.680 96.030 104.855 ;
        RECT 89.255 104.390 91.410 104.670 ;
        RECT 86.460 104.265 86.790 104.370 ;
        RECT 85.320 104.095 86.290 104.200 ;
        RECT 87.025 104.095 87.370 104.200 ;
        RECT 85.320 103.925 87.370 104.095 ;
        RECT 87.700 103.755 87.870 104.390 ;
        RECT 90.420 104.355 91.410 104.390 ;
        RECT 88.040 103.860 88.670 104.215 ;
        RECT 84.980 103.585 86.330 103.755 ;
        RECT 86.785 103.690 87.870 103.755 ;
        RECT 86.785 103.585 88.330 103.690 ;
        RECT 81.860 102.535 82.430 102.865 ;
        RECT 81.520 102.110 82.040 102.365 ;
        RECT 79.880 101.860 80.210 101.885 ;
        RECT 79.880 101.690 80.220 101.860 ;
        RECT 80.390 101.715 81.620 101.885 ;
        RECT 82.260 101.860 82.430 102.535 ;
        RECT 82.600 102.980 82.940 103.290 ;
        RECT 83.110 102.980 83.745 103.295 ;
        RECT 84.980 103.290 85.150 103.585 ;
        RECT 87.700 103.520 88.330 103.585 ;
        RECT 87.700 103.295 87.870 103.520 ;
        RECT 88.500 103.350 88.670 103.860 ;
        RECT 83.915 103.250 85.150 103.290 ;
        RECT 83.915 103.000 85.610 103.250 ;
        RECT 85.780 103.040 87.070 103.295 ;
        RECT 87.240 103.040 87.870 103.295 ;
        RECT 83.915 102.980 85.150 103.000 ;
        RECT 82.600 102.430 82.770 102.980 ;
        RECT 82.940 102.600 84.810 102.810 ;
        RECT 84.130 102.575 84.810 102.600 ;
        RECT 82.600 102.100 83.230 102.430 ;
        RECT 83.790 102.260 83.960 102.320 ;
        RECT 82.260 101.815 82.890 101.860 ;
        RECT 79.880 101.605 80.210 101.690 ;
        RECT 79.105 101.185 80.210 101.435 ;
        RECT 79.105 100.815 79.710 101.185 ;
        RECT 77.855 100.465 79.710 100.815 ;
        RECT 79.105 99.235 79.710 100.465 ;
        RECT 79.880 100.940 80.210 101.015 ;
        RECT 79.880 100.770 80.220 100.940 ;
        RECT 79.880 100.765 80.210 100.770 ;
        RECT 79.880 100.175 80.050 100.765 ;
        RECT 80.390 100.595 80.560 101.715 ;
        RECT 81.440 101.475 81.620 101.715 ;
        RECT 81.790 101.690 82.890 101.815 ;
        RECT 81.790 101.645 82.430 101.690 ;
        RECT 81.070 101.300 81.270 101.460 ;
        RECT 80.220 100.345 80.560 100.595 ;
        RECT 79.880 99.925 80.210 100.175 ;
        RECT 80.390 99.955 80.560 100.345 ;
        RECT 80.730 101.130 81.270 101.300 ;
        RECT 81.440 101.145 82.090 101.475 ;
        RECT 80.730 100.295 80.900 101.130 ;
        RECT 81.070 100.465 81.270 100.960 ;
        RECT 81.440 100.635 81.620 101.145 ;
        RECT 82.260 100.975 82.430 101.645 ;
        RECT 83.060 101.460 83.230 102.100 ;
        RECT 83.420 101.765 83.960 102.260 ;
        RECT 82.600 101.130 83.230 101.460 ;
        RECT 81.790 100.950 82.430 100.975 ;
        RECT 81.790 100.805 82.890 100.950 ;
        RECT 82.260 100.780 82.890 100.805 ;
        RECT 81.440 100.305 82.090 100.635 ;
        RECT 80.730 100.125 81.270 100.295 ;
        RECT 82.260 100.135 82.430 100.780 ;
        RECT 83.060 100.600 83.230 101.130 ;
        RECT 83.420 100.785 83.620 101.585 ;
        RECT 83.790 100.615 83.960 101.765 ;
        RECT 84.130 101.460 84.310 102.575 ;
        RECT 84.980 102.450 85.150 102.980 ;
        RECT 85.780 102.790 85.950 103.040 ;
        RECT 85.320 102.620 85.950 102.790 ;
        RECT 86.120 102.660 86.710 102.830 ;
        RECT 84.980 102.405 85.950 102.450 ;
        RECT 84.520 102.200 85.950 102.405 ;
        RECT 84.520 102.075 85.150 102.200 ;
        RECT 84.480 101.690 84.810 101.880 ;
        RECT 84.130 101.160 84.470 101.460 ;
        RECT 84.640 100.990 84.810 101.690 ;
        RECT 84.130 100.770 84.810 100.990 ;
        RECT 84.980 101.570 85.150 102.075 ;
        RECT 85.360 101.780 85.950 102.030 ;
        RECT 84.980 101.240 85.610 101.570 ;
        RECT 82.600 100.270 83.230 100.600 ;
        RECT 83.400 100.285 83.960 100.615 ;
        RECT 84.980 100.600 85.150 101.240 ;
        RECT 85.780 101.050 85.950 101.780 ;
        RECT 85.360 100.800 85.950 101.050 ;
        RECT 85.780 100.740 85.950 100.800 ;
        RECT 86.120 100.850 86.290 102.660 ;
        RECT 86.540 102.500 86.710 102.660 ;
        RECT 86.900 102.790 87.070 103.040 ;
        RECT 87.700 102.850 87.870 103.040 ;
        RECT 88.040 103.020 88.670 103.350 ;
        RECT 88.840 103.065 89.110 104.215 ;
        RECT 89.280 103.860 90.250 104.215 ;
        RECT 89.280 103.350 89.450 103.860 ;
        RECT 90.420 103.690 90.590 104.355 ;
        RECT 91.580 104.325 92.150 104.670 ;
        RECT 92.320 104.340 92.905 104.670 ;
        RECT 93.140 104.390 94.035 104.680 ;
        RECT 94.695 104.390 96.030 104.680 ;
        RECT 90.930 104.150 91.100 104.160 ;
        RECT 90.800 103.980 92.150 104.150 ;
        RECT 89.620 103.520 90.590 103.690 ;
        RECT 86.900 102.620 87.530 102.790 ;
        RECT 87.700 102.430 88.330 102.850 ;
        RECT 87.320 102.370 88.330 102.430 ;
        RECT 87.240 102.340 88.330 102.370 ;
        RECT 86.460 102.115 87.025 102.320 ;
        RECT 87.240 102.200 87.870 102.340 ;
        RECT 86.460 101.990 86.790 102.115 ;
        RECT 87.320 102.100 87.870 102.200 ;
        RECT 88.500 102.130 88.670 103.020 ;
        RECT 89.280 103.020 90.250 103.350 ;
        RECT 90.420 103.190 90.590 103.520 ;
        RECT 90.800 103.460 91.730 103.810 ;
        RECT 91.900 103.595 92.150 103.980 ;
        RECT 92.320 103.810 92.500 104.340 ;
        RECT 93.140 104.170 93.310 104.390 ;
        RECT 92.670 104.000 93.310 104.170 ;
        RECT 92.320 103.580 92.905 103.810 ;
        RECT 91.170 103.425 91.730 103.460 ;
        RECT 91.170 103.405 92.150 103.425 ;
        RECT 91.170 103.255 92.905 103.405 ;
        RECT 87.190 101.855 87.360 101.860 ;
        RECT 86.920 101.760 87.385 101.855 ;
        RECT 86.525 101.685 87.385 101.760 ;
        RECT 86.525 101.590 87.090 101.685 ;
        RECT 87.700 101.630 87.870 102.100 ;
        RECT 88.040 101.800 88.670 102.130 ;
        RECT 88.840 102.085 89.110 102.895 ;
        RECT 89.280 102.510 89.450 103.020 ;
        RECT 89.620 102.680 90.250 102.850 ;
        RECT 89.280 102.180 89.910 102.510 ;
        RECT 86.540 101.430 86.710 101.590 ;
        RECT 86.915 101.210 87.370 101.420 ;
        RECT 87.700 101.300 88.330 101.630 ;
        RECT 86.915 101.200 87.085 101.210 ;
        RECT 86.460 101.030 87.085 101.200 ;
        RECT 87.280 100.925 87.450 101.010 ;
        RECT 87.280 100.850 87.530 100.925 ;
        RECT 84.130 100.270 85.150 100.600 ;
        RECT 86.120 100.680 87.530 100.850 ;
        RECT 86.120 100.510 86.290 100.680 ;
        RECT 87.700 100.510 87.870 101.300 ;
        RECT 88.500 101.130 88.670 101.800 ;
        RECT 85.320 100.340 86.290 100.510 ;
        RECT 86.460 100.295 87.030 100.490 ;
        RECT 80.390 99.785 80.900 99.955 ;
        RECT 79.880 99.615 80.220 99.720 ;
        RECT 79.880 99.405 80.560 99.615 ;
        RECT 79.105 98.985 80.210 99.235 ;
        RECT 79.105 98.875 79.710 98.985 ;
        RECT 76.275 98.700 76.990 98.875 ;
        RECT 79.540 98.700 79.710 98.875 ;
        RECT 80.390 98.815 80.560 99.405 ;
        RECT 76.275 97.955 77.535 98.700 ;
        RECT 72.540 96.730 72.710 97.220 ;
        RECT 73.250 97.150 73.930 97.920 ;
        RECT 72.880 96.730 73.590 96.980 ;
        RECT 71.020 96.520 71.550 96.565 ;
        RECT 72.190 96.520 72.370 96.690 ;
        RECT 72.880 96.520 73.090 96.730 ;
        RECT 73.760 96.560 73.930 97.150 ;
        RECT 71.020 96.350 72.020 96.520 ;
        RECT 71.020 96.235 71.550 96.350 ;
        RECT 70.680 96.010 71.210 96.030 ;
        RECT 69.350 95.710 71.210 96.010 ;
        RECT 71.380 95.850 71.550 96.235 ;
        RECT 72.190 96.110 73.090 96.520 ;
        RECT 73.260 96.310 73.930 96.560 ;
        RECT 74.100 97.780 74.270 97.955 ;
        RECT 76.820 97.780 77.535 97.955 ;
        RECT 74.100 95.850 74.705 97.780 ;
        RECT 76.275 97.115 77.535 97.780 ;
        RECT 79.105 98.395 79.710 98.700 ;
        RECT 79.880 98.565 80.560 98.815 ;
        RECT 79.105 98.090 80.210 98.395 ;
        RECT 76.275 96.775 78.365 97.115 ;
        RECT 76.275 96.195 77.535 96.775 ;
        RECT 75.445 95.855 77.535 96.195 ;
        RECT 71.380 95.550 72.030 95.850 ;
        RECT 69.000 95.235 69.670 95.540 ;
        RECT 71.380 95.530 71.550 95.550 ;
        RECT 69.840 95.250 70.470 95.525 ;
        RECT 70.640 95.200 71.550 95.530 ;
        RECT 72.200 95.410 73.185 95.850 ;
        RECT 73.355 95.580 74.705 95.850 ;
        RECT 72.200 95.380 73.925 95.410 ;
        RECT 64.650 94.960 66.770 95.020 ;
        RECT 62.130 94.270 65.020 94.790 ;
        RECT 65.190 94.745 66.770 94.960 ;
        RECT 65.190 94.270 66.110 94.745 ;
        RECT 66.950 94.590 67.470 95.020 ;
        RECT 67.650 94.760 68.830 95.020 ;
        RECT 66.950 94.575 68.490 94.590 ;
        RECT 66.280 94.420 68.490 94.575 ;
        RECT 66.280 94.405 67.470 94.420 ;
        RECT 66.280 94.325 66.740 94.405 ;
        RECT 67.820 94.315 68.490 94.420 ;
        RECT 62.130 93.995 63.390 94.270 ;
        RECT 65.940 94.150 66.110 94.270 ;
        RECT 60.500 91.970 61.440 93.830 ;
        RECT 62.130 93.825 63.850 93.995 ;
        RECT 62.130 93.660 63.390 93.825 ;
        RECT 61.610 93.155 63.390 93.660 ;
        RECT 64.020 93.670 65.370 94.100 ;
        RECT 65.940 94.075 66.605 94.150 ;
        RECT 65.540 93.820 66.605 94.075 ;
        RECT 67.020 94.005 67.620 94.235 ;
        RECT 68.660 94.115 68.830 94.760 ;
        RECT 65.540 93.745 66.110 93.820 ;
        RECT 64.020 93.655 64.190 93.670 ;
        RECT 63.560 93.325 64.190 93.655 ;
        RECT 65.200 93.575 65.370 93.670 ;
        RECT 64.360 93.330 65.030 93.500 ;
        RECT 65.200 93.405 65.640 93.575 ;
        RECT 61.610 92.985 64.190 93.155 ;
        RECT 61.610 91.970 63.390 92.985 ;
        RECT 64.360 92.580 64.530 93.330 ;
        RECT 65.940 93.235 66.110 93.745 ;
        RECT 66.775 93.640 67.270 93.820 ;
        RECT 66.330 93.410 67.270 93.640 ;
        RECT 67.450 93.675 67.620 94.005 ;
        RECT 67.815 93.900 68.830 94.115 ;
        RECT 67.450 93.425 67.915 93.675 ;
        RECT 67.450 93.240 67.620 93.425 ;
        RECT 68.150 93.240 68.490 93.715 ;
        RECT 68.660 93.655 68.830 93.900 ;
        RECT 69.050 93.825 69.340 95.020 ;
        RECT 69.510 94.670 69.970 95.000 ;
        RECT 70.140 94.670 70.470 95.020 ;
        RECT 70.640 94.745 71.160 95.000 ;
        RECT 71.380 94.950 71.550 95.200 ;
        RECT 71.745 95.120 73.925 95.380 ;
        RECT 69.510 94.005 69.680 94.670 ;
        RECT 69.850 94.275 70.470 94.500 ;
        RECT 69.510 93.835 69.970 94.005 ;
        RECT 68.660 93.375 69.630 93.655 ;
        RECT 69.800 93.505 69.970 93.835 ;
        RECT 70.140 93.675 70.470 94.275 ;
        RECT 70.640 94.075 70.810 94.745 ;
        RECT 71.380 94.690 72.030 94.950 ;
        RECT 71.380 94.575 71.550 94.690 ;
        RECT 70.980 94.245 71.550 94.575 ;
        RECT 72.200 94.685 73.185 95.120 ;
        RECT 74.100 94.950 74.705 95.580 ;
        RECT 73.370 94.695 74.705 94.950 ;
        RECT 72.200 94.510 72.370 94.685 ;
        RECT 71.745 94.250 72.370 94.510 ;
        RECT 71.380 94.080 71.550 94.245 ;
        RECT 70.640 93.905 71.160 94.075 ;
        RECT 70.640 93.505 70.810 93.905 ;
        RECT 71.380 93.830 72.030 94.080 ;
        RECT 71.380 93.735 71.550 93.830 ;
        RECT 64.700 92.750 65.260 93.160 ;
        RECT 65.430 92.920 66.110 93.235 ;
        RECT 65.430 92.580 65.770 92.690 ;
        RECT 64.360 92.400 65.770 92.580 ;
        RECT 64.185 92.040 64.530 92.400 ;
        RECT 65.940 92.260 66.110 92.920 ;
        RECT 66.330 92.985 67.620 93.240 ;
        RECT 66.330 92.450 66.595 92.985 ;
        RECT 66.790 92.430 67.270 92.815 ;
        RECT 67.450 92.700 67.620 92.985 ;
        RECT 67.790 93.060 67.980 93.200 ;
        RECT 68.660 93.060 68.830 93.375 ;
        RECT 69.800 93.335 70.810 93.505 ;
        RECT 70.980 93.355 71.550 93.735 ;
        RECT 72.200 93.650 72.370 94.250 ;
        RECT 71.745 93.390 72.370 93.650 ;
        RECT 70.140 93.230 70.470 93.335 ;
        RECT 71.380 93.220 71.550 93.355 ;
        RECT 67.790 92.870 68.830 93.060 ;
        RECT 69.000 93.060 69.970 93.165 ;
        RECT 70.705 93.060 71.050 93.165 ;
        RECT 69.000 92.890 71.050 93.060 ;
        RECT 71.380 92.970 72.030 93.220 ;
        RECT 68.155 92.720 68.830 92.870 ;
        RECT 71.380 92.720 71.550 92.970 ;
        RECT 72.200 92.790 72.370 93.390 ;
        RECT 67.450 92.445 67.985 92.700 ;
        RECT 68.155 92.430 70.035 92.720 ;
        RECT 70.550 92.430 71.550 92.720 ;
        RECT 71.745 92.530 72.370 92.790 ;
        RECT 68.660 92.260 68.830 92.430 ;
        RECT 65.940 92.230 66.910 92.260 ;
        RECT 64.700 92.035 65.260 92.230 ;
        RECT 65.090 92.030 65.260 92.035 ;
        RECT 65.430 91.990 66.910 92.230 ;
        RECT 60.500 91.800 60.670 91.970 ;
        RECT 63.220 91.800 63.390 91.970 ;
        RECT 65.940 91.880 66.910 91.990 ;
        RECT 65.940 91.800 66.110 91.880 ;
        RECT 60.500 91.510 61.395 91.800 ;
        RECT 62.055 91.510 64.555 91.800 ;
        RECT 65.215 91.510 66.110 91.800 ;
        RECT 60.500 89.890 60.670 91.510 ;
        RECT 63.220 91.340 63.390 91.510 ;
        RECT 65.940 91.340 66.110 91.510 ;
        RECT 60.840 90.900 61.070 91.230 ;
        RECT 61.240 91.060 62.250 91.340 ;
        RECT 63.220 91.235 64.480 91.340 ;
        RECT 60.840 90.310 61.050 90.900 ;
        RECT 61.240 90.480 61.490 91.060 ;
        RECT 60.840 90.060 61.470 90.310 ;
        RECT 61.660 90.140 61.910 90.890 ;
        RECT 62.080 90.810 62.250 91.060 ;
        RECT 62.420 90.980 64.480 91.235 ;
        RECT 62.080 90.480 63.050 90.810 ;
        RECT 60.500 89.720 61.130 89.890 ;
        RECT 60.500 89.040 60.670 89.720 ;
        RECT 61.300 89.550 61.470 90.060 ;
        RECT 62.080 89.970 62.250 90.480 ;
        RECT 63.220 90.420 64.480 90.980 ;
        RECT 64.650 91.290 66.110 91.340 ;
        RECT 64.650 90.960 66.490 91.290 ;
        RECT 64.650 90.590 66.110 90.960 ;
        RECT 63.220 90.310 65.000 90.420 ;
        RECT 62.420 90.140 65.000 90.310 ;
        RECT 60.840 89.210 61.470 89.550 ;
        RECT 61.660 89.210 61.910 89.970 ;
        RECT 62.080 89.640 63.050 89.970 ;
        RECT 63.220 89.670 65.000 90.140 ;
        RECT 65.170 89.670 66.110 90.590 ;
        RECT 63.220 89.470 63.390 89.670 ;
        RECT 62.080 89.210 63.390 89.470 ;
        RECT 63.560 89.240 64.230 89.410 ;
        RECT 63.220 89.070 63.390 89.210 ;
        RECT 63.220 89.040 63.890 89.070 ;
        RECT 60.500 87.455 61.215 89.040 ;
        RECT 62.785 88.740 63.890 89.040 ;
        RECT 64.060 88.975 64.230 89.240 ;
        RECT 64.400 89.145 65.050 89.495 ;
        RECT 65.220 89.240 65.680 89.410 ;
        RECT 65.220 88.975 65.390 89.240 ;
        RECT 65.940 89.070 66.110 89.670 ;
        RECT 64.060 88.745 65.390 88.975 ;
        RECT 65.560 88.740 66.110 89.070 ;
        RECT 66.320 89.010 66.490 90.770 ;
        RECT 66.660 90.020 66.930 91.710 ;
        RECT 67.100 91.135 67.300 92.260 ;
        RECT 67.470 91.880 68.830 92.260 ;
        RECT 68.660 91.800 68.830 91.880 ;
        RECT 71.380 92.360 71.550 92.430 ;
        RECT 71.380 92.115 72.030 92.360 ;
        RECT 71.380 91.800 71.550 92.115 ;
        RECT 72.200 91.945 72.370 92.530 ;
        RECT 67.130 91.110 67.300 91.135 ;
        RECT 67.470 91.380 68.490 91.710 ;
        RECT 68.660 91.510 69.995 91.800 ;
        RECT 70.655 91.510 71.550 91.800 ;
        RECT 71.745 91.670 72.370 91.945 ;
        RECT 67.100 89.735 67.300 90.825 ;
        RECT 67.470 90.350 67.690 91.380 ;
        RECT 68.660 91.340 68.830 91.510 ;
        RECT 71.380 91.500 71.550 91.510 ;
        RECT 71.380 91.340 72.030 91.500 ;
        RECT 68.660 91.210 69.920 91.340 ;
        RECT 67.860 90.650 69.920 91.210 ;
        RECT 70.090 91.255 72.030 91.340 ;
        RECT 70.090 90.820 71.550 91.255 ;
        RECT 72.200 91.085 72.370 91.670 ;
        RECT 71.745 90.825 72.370 91.085 ;
        RECT 70.630 90.655 71.550 90.820 ;
        RECT 67.860 90.520 70.460 90.650 ;
        RECT 67.470 90.020 68.490 90.350 ;
        RECT 68.660 90.130 70.460 90.520 ;
        RECT 70.630 90.395 72.030 90.655 ;
        RECT 70.630 90.130 71.550 90.395 ;
        RECT 72.200 90.225 72.370 90.825 ;
        RECT 67.470 89.510 67.690 90.020 ;
        RECT 68.660 89.850 68.830 90.130 ;
        RECT 67.860 89.680 68.830 89.850 ;
        RECT 69.000 89.700 69.670 89.870 ;
        RECT 68.660 89.530 68.830 89.680 ;
        RECT 66.660 89.180 68.490 89.510 ;
        RECT 68.660 89.200 69.330 89.530 ;
        RECT 69.500 89.435 69.670 89.700 ;
        RECT 69.840 89.605 70.490 89.955 ;
        RECT 70.660 89.700 71.120 89.870 ;
        RECT 71.380 89.795 71.550 90.130 ;
        RECT 71.745 89.965 72.370 90.225 ;
        RECT 70.660 89.435 70.830 89.700 ;
        RECT 71.380 89.535 72.030 89.795 ;
        RECT 71.380 89.530 71.550 89.535 ;
        RECT 69.500 89.205 70.830 89.435 ;
        RECT 71.000 89.200 71.550 89.530 ;
        RECT 72.200 89.365 72.370 89.965 ;
        RECT 68.660 89.010 68.830 89.200 ;
        RECT 66.320 88.755 66.810 89.010 ;
        RECT 67.020 88.755 67.350 88.995 ;
        RECT 67.520 88.755 68.830 89.010 ;
        RECT 69.000 88.845 71.120 89.030 ;
        RECT 71.380 88.935 71.550 89.200 ;
        RECT 71.745 89.105 72.370 89.365 ;
        RECT 62.785 88.145 63.390 88.740 ;
        RECT 65.940 88.580 66.110 88.740 ;
        RECT 68.660 88.605 68.830 88.755 ;
        RECT 71.380 88.675 72.110 88.935 ;
        RECT 63.560 88.385 65.680 88.570 ;
        RECT 65.940 88.250 66.590 88.580 ;
        RECT 66.775 88.255 67.350 88.570 ;
        RECT 67.695 88.300 68.490 88.520 ;
        RECT 68.660 88.340 69.290 88.605 ;
        RECT 69.800 88.395 70.750 88.675 ;
        RECT 71.380 88.590 71.550 88.675 ;
        RECT 70.920 88.340 71.550 88.590 ;
        RECT 72.540 88.505 72.790 94.515 ;
        RECT 72.960 94.510 73.185 94.685 ;
        RECT 72.960 94.250 73.925 94.510 ;
        RECT 74.095 94.375 74.705 94.695 ;
        RECT 72.960 93.650 73.200 94.250 ;
        RECT 74.095 94.080 75.955 94.375 ;
        RECT 73.370 94.025 75.955 94.080 ;
        RECT 73.370 93.835 74.705 94.025 ;
        RECT 72.960 93.390 73.925 93.650 ;
        RECT 72.960 92.790 73.200 93.390 ;
        RECT 74.095 93.220 74.705 93.835 ;
        RECT 73.370 92.975 74.705 93.220 ;
        RECT 72.960 92.530 73.925 92.790 ;
        RECT 72.960 91.945 73.200 92.530 ;
        RECT 74.095 92.435 74.705 92.975 ;
        RECT 76.275 93.355 77.535 95.855 ;
        RECT 79.105 95.940 79.710 98.090 ;
        RECT 80.390 97.920 80.560 98.565 ;
        RECT 79.880 97.150 80.560 97.920 ;
        RECT 80.730 97.390 80.900 99.785 ;
        RECT 81.070 98.775 81.270 100.125 ;
        RECT 81.790 100.080 82.430 100.135 ;
        RECT 84.980 100.080 85.150 100.270 ;
        RECT 87.220 100.250 87.870 100.510 ;
        RECT 81.790 99.965 83.720 100.080 ;
        RECT 81.440 99.365 82.090 99.695 ;
        RECT 82.260 99.560 83.720 99.965 ;
        RECT 83.890 99.625 85.150 100.080 ;
        RECT 87.700 100.065 87.870 100.250 ;
        RECT 85.320 99.795 85.930 100.055 ;
        RECT 81.440 98.855 81.620 99.365 ;
        RECT 82.260 99.195 83.180 99.560 ;
        RECT 83.890 99.390 85.510 99.625 ;
        RECT 81.790 99.025 83.180 99.195 ;
        RECT 82.260 98.870 83.180 99.025 ;
        RECT 83.350 99.295 85.510 99.390 ;
        RECT 83.350 98.870 85.150 99.295 ;
        RECT 85.680 99.115 85.930 99.795 ;
        RECT 85.320 98.945 85.930 99.115 ;
        RECT 81.440 98.605 82.090 98.855 ;
        RECT 81.070 97.915 81.270 98.585 ;
        RECT 81.440 98.050 81.700 98.380 ;
        RECT 80.730 97.220 81.270 97.390 ;
        RECT 79.880 96.560 80.050 97.150 ;
        RECT 80.220 96.730 80.930 96.980 ;
        RECT 81.100 96.730 81.270 97.220 ;
        RECT 81.440 97.020 81.620 98.050 ;
        RECT 81.870 97.625 82.090 98.605 ;
        RECT 82.260 98.700 82.430 98.870 ;
        RECT 84.980 98.700 85.150 98.870 ;
        RECT 82.260 98.350 83.230 98.700 ;
        RECT 83.980 98.690 85.150 98.700 ;
        RECT 83.980 98.520 85.590 98.690 ;
        RECT 83.980 98.350 85.150 98.520 ;
        RECT 85.760 98.350 85.930 98.945 ;
        RECT 82.260 97.720 82.430 98.350 ;
        RECT 82.600 97.890 84.735 98.180 ;
        RECT 84.980 97.720 85.150 98.350 ;
        RECT 82.260 97.460 83.210 97.720 ;
        RECT 82.260 97.360 82.790 97.460 ;
        RECT 81.790 97.190 82.790 97.360 ;
        RECT 83.420 97.290 83.670 97.720 ;
        RECT 83.840 97.470 85.150 97.720 ;
        RECT 79.880 96.310 80.550 96.560 ;
        RECT 80.720 96.520 80.930 96.730 ;
        RECT 81.440 96.690 81.700 97.020 ;
        RECT 82.260 96.775 82.790 97.190 ;
        RECT 82.960 97.080 84.810 97.290 ;
        RECT 81.440 96.520 81.620 96.690 ;
        RECT 82.260 96.520 82.430 96.775 ;
        RECT 82.960 96.605 83.130 97.080 ;
        RECT 83.840 97.000 84.810 97.080 ;
        RECT 80.720 96.110 81.620 96.520 ;
        RECT 81.790 96.350 82.430 96.520 ;
        RECT 82.600 96.365 83.130 96.605 ;
        RECT 83.340 96.825 83.670 96.900 ;
        RECT 83.340 96.530 84.700 96.825 ;
        RECT 82.260 96.195 82.430 96.350 ;
        RECT 82.260 95.940 82.790 96.195 ;
        RECT 79.105 95.680 80.720 95.940 ;
        RECT 79.105 95.295 79.710 95.680 ;
        RECT 80.900 95.510 81.420 95.940 ;
        RECT 81.600 95.865 82.790 95.940 ;
        RECT 81.600 95.665 82.430 95.865 ;
        RECT 82.960 95.695 83.130 96.365 ;
        RECT 83.340 96.050 84.700 96.360 ;
        RECT 77.855 95.035 79.710 95.295 ;
        RECT 79.880 95.495 81.420 95.510 ;
        RECT 79.880 95.340 82.090 95.495 ;
        RECT 79.880 95.235 80.550 95.340 ;
        RECT 80.900 95.325 82.090 95.340 ;
        RECT 81.630 95.245 82.090 95.325 ;
        RECT 77.855 94.945 80.555 95.035 ;
        RECT 79.105 94.820 80.555 94.945 ;
        RECT 80.750 94.925 81.350 95.155 ;
        RECT 82.260 95.070 82.430 95.665 ;
        RECT 82.600 95.450 83.130 95.695 ;
        RECT 83.340 95.590 84.085 95.880 ;
        RECT 83.300 95.280 84.085 95.420 ;
        RECT 79.105 93.980 79.710 94.820 ;
        RECT 79.880 94.160 80.220 94.635 ;
        RECT 80.750 94.595 80.920 94.925 ;
        RECT 81.765 94.740 82.430 95.070 ;
        RECT 82.635 95.010 84.085 95.280 ;
        RECT 84.260 95.385 84.810 95.715 ;
        RECT 82.635 94.790 83.170 95.010 ;
        RECT 80.455 94.345 80.920 94.595 ;
        RECT 80.750 94.160 80.920 94.345 ;
        RECT 81.100 94.560 81.595 94.740 ;
        RECT 82.260 94.620 82.430 94.740 ;
        RECT 81.100 94.330 82.040 94.560 ;
        RECT 82.260 94.270 83.150 94.620 ;
        RECT 83.340 94.270 84.085 94.840 ;
        RECT 84.260 94.695 84.430 95.385 ;
        RECT 84.980 95.195 85.150 97.470 ;
        RECT 85.320 98.020 85.930 98.350 ;
        RECT 86.110 99.520 86.750 100.020 ;
        RECT 86.920 99.770 87.870 100.065 ;
        RECT 88.040 100.800 88.670 101.130 ;
        RECT 88.840 101.100 89.110 101.915 ;
        RECT 89.280 101.640 89.910 101.970 ;
        RECT 89.280 101.130 89.450 101.640 ;
        RECT 90.080 101.470 90.250 102.680 ;
        RECT 89.620 101.300 90.250 101.470 ;
        RECT 90.420 102.785 90.990 103.190 ;
        RECT 90.420 101.915 90.590 102.785 ;
        RECT 90.420 101.585 90.990 101.915 ;
        RECT 91.170 101.895 91.340 103.255 ;
        RECT 91.980 103.235 92.905 103.255 ;
        RECT 92.535 103.160 92.905 103.235 ;
        RECT 91.510 102.990 91.870 103.085 ;
        RECT 91.510 102.820 92.830 102.990 ;
        RECT 91.510 102.065 91.730 102.820 ;
        RECT 92.125 102.645 92.455 102.650 ;
        RECT 92.125 102.480 92.490 102.645 ;
        RECT 92.660 102.530 92.830 102.820 ;
        RECT 93.140 102.855 93.310 104.000 ;
        RECT 95.860 103.740 96.030 104.390 ;
        RECT 98.580 104.850 99.520 104.855 ;
        RECT 99.690 104.850 101.470 105.600 ;
        RECT 104.020 105.540 105.480 105.940 ;
        RECT 105.650 105.950 107.825 106.060 ;
        RECT 105.650 105.600 106.910 105.950 ;
        RECT 108.945 105.940 110.175 106.110 ;
        RECT 109.460 105.600 110.175 105.940 ;
        RECT 104.020 105.120 104.940 105.540 ;
        RECT 105.650 105.370 108.000 105.600 ;
        RECT 102.830 105.075 103.000 105.080 ;
        RECT 98.580 104.680 98.750 104.850 ;
        RECT 101.300 104.680 101.470 104.850 ;
        RECT 102.265 104.710 102.610 105.070 ;
        RECT 102.780 104.880 103.340 105.075 ;
        RECT 103.510 104.880 104.940 105.120 ;
        RECT 104.020 104.850 104.940 104.880 ;
        RECT 105.110 104.910 108.000 105.370 ;
        RECT 108.170 105.315 110.175 105.600 ;
        RECT 111.745 105.315 112.350 106.905 ;
        RECT 108.170 105.080 109.630 105.315 ;
        RECT 105.110 104.850 108.540 104.910 ;
        RECT 98.580 104.390 99.475 104.680 ;
        RECT 100.135 104.390 101.470 104.680 ;
        RECT 98.580 103.755 98.750 104.390 ;
        RECT 101.300 104.125 101.470 104.390 ;
        RECT 102.440 104.530 103.850 104.710 ;
        RECT 101.300 103.955 102.270 104.125 ;
        RECT 95.860 103.410 96.880 103.740 ;
        RECT 93.530 103.025 94.050 103.280 ;
        RECT 92.320 102.360 92.490 102.480 ;
        RECT 93.140 102.525 93.710 102.855 ;
        RECT 91.170 101.725 91.780 101.895 ;
        RECT 91.950 101.840 92.150 102.310 ;
        RECT 92.320 102.140 92.845 102.360 ;
        RECT 93.140 102.015 93.310 102.525 ;
        RECT 93.880 102.355 94.050 103.025 ;
        RECT 94.220 102.950 94.550 103.300 ;
        RECT 94.720 102.950 95.180 103.280 ;
        RECT 93.530 102.185 94.050 102.355 ;
        RECT 93.140 101.860 93.710 102.015 ;
        RECT 91.610 101.670 91.780 101.725 ;
        RECT 92.475 101.690 93.710 101.860 ;
        RECT 89.280 100.800 90.250 101.130 ;
        RECT 90.420 100.990 90.590 101.585 ;
        RECT 91.610 101.500 92.230 101.670 ;
        RECT 93.140 101.635 93.710 101.690 ;
        RECT 93.880 101.785 94.050 102.185 ;
        RECT 94.220 102.555 94.840 102.780 ;
        RECT 94.220 101.955 94.550 102.555 ;
        RECT 95.010 102.285 95.180 102.950 ;
        RECT 94.720 102.115 95.180 102.285 ;
        RECT 94.720 101.785 94.890 102.115 ;
        RECT 95.350 102.105 95.640 103.300 ;
        RECT 95.860 101.935 96.030 103.410 ;
        RECT 97.050 103.395 97.610 103.725 ;
        RECT 97.780 103.410 98.410 103.740 ;
        RECT 98.580 103.420 99.250 103.755 ;
        RECT 96.200 103.020 96.880 103.240 ;
        RECT 96.200 102.320 96.370 103.020 ;
        RECT 96.540 102.550 96.880 102.850 ;
        RECT 96.200 102.130 96.530 102.320 ;
        RECT 90.760 101.400 91.430 101.415 ;
        RECT 90.760 101.330 91.440 101.400 ;
        RECT 92.400 101.330 92.970 101.495 ;
        RECT 90.760 101.160 92.970 101.330 ;
        RECT 93.140 101.000 93.310 101.635 ;
        RECT 93.880 101.615 94.890 101.785 ;
        RECT 95.060 101.655 96.490 101.935 ;
        RECT 94.220 101.510 94.550 101.615 ;
        RECT 95.860 101.605 96.490 101.655 ;
        RECT 93.640 101.340 93.985 101.445 ;
        RECT 94.720 101.340 95.690 101.445 ;
        RECT 93.640 101.170 95.690 101.340 ;
        RECT 95.860 101.030 96.030 101.605 ;
        RECT 96.700 101.435 96.880 102.550 ;
        RECT 97.050 102.245 97.220 103.395 ;
        RECT 97.390 102.425 97.590 103.225 ;
        RECT 97.780 102.880 97.950 103.410 ;
        RECT 98.580 103.230 98.750 103.420 ;
        RECT 99.420 103.405 99.990 103.760 ;
        RECT 100.160 103.435 100.620 103.760 ;
        RECT 100.110 103.235 100.280 103.240 ;
        RECT 98.120 103.060 98.750 103.230 ;
        RECT 97.780 102.550 98.410 102.880 ;
        RECT 98.580 102.850 98.750 103.060 ;
        RECT 98.970 103.050 99.490 103.220 ;
        RECT 97.050 101.750 97.590 102.245 ;
        RECT 97.780 101.910 97.950 102.550 ;
        RECT 98.580 102.520 99.150 102.850 ;
        RECT 98.580 102.320 98.750 102.520 ;
        RECT 99.320 102.350 99.490 103.050 ;
        RECT 99.660 102.525 100.280 103.235 ;
        RECT 98.120 102.150 98.750 102.320 ;
        RECT 98.970 102.180 99.490 102.350 ;
        RECT 98.580 102.010 98.750 102.150 ;
        RECT 97.780 101.580 98.410 101.910 ;
        RECT 96.200 101.410 96.880 101.435 ;
        RECT 96.200 101.200 98.070 101.410 ;
        RECT 98.240 101.030 98.410 101.580 ;
        RECT 95.860 101.000 97.095 101.030 ;
        RECT 93.140 100.990 94.140 101.000 ;
        RECT 88.040 100.130 88.210 100.800 ;
        RECT 89.280 100.630 89.450 100.800 ;
        RECT 90.420 100.735 91.815 100.990 ;
        RECT 92.315 100.735 94.140 100.990 ;
        RECT 90.420 100.630 90.590 100.735 ;
        RECT 88.380 100.300 89.450 100.630 ;
        RECT 89.620 100.540 90.590 100.630 ;
        RECT 93.140 100.710 94.140 100.735 ;
        RECT 94.655 100.720 97.095 101.000 ;
        RECT 94.655 100.710 96.030 100.720 ;
        RECT 97.265 100.715 97.900 101.030 ;
        RECT 98.070 100.720 98.410 101.030 ;
        RECT 98.580 101.630 99.150 102.010 ;
        RECT 99.320 101.780 99.490 102.180 ;
        RECT 99.660 101.950 99.990 102.355 ;
        RECT 100.450 102.335 100.620 103.435 ;
        RECT 100.160 102.165 100.620 102.335 ;
        RECT 100.160 101.780 100.330 102.165 ;
        RECT 100.790 102.100 101.080 103.760 ;
        RECT 101.300 103.285 101.470 103.955 ;
        RECT 101.640 103.455 102.270 103.785 ;
        RECT 102.440 103.780 102.610 104.530 ;
        RECT 103.510 104.420 103.850 104.530 ;
        RECT 104.020 104.680 104.190 104.850 ;
        RECT 106.740 104.680 108.540 104.850 ;
        RECT 104.020 104.390 104.915 104.680 ;
        RECT 105.575 104.390 108.540 104.680 ;
        RECT 108.710 104.680 109.630 105.080 ;
        RECT 112.180 104.680 112.350 105.315 ;
        RECT 108.710 104.390 110.355 104.680 ;
        RECT 111.015 104.390 112.350 104.680 ;
        RECT 102.780 103.950 103.340 104.360 ;
        RECT 104.020 104.220 104.190 104.390 ;
        RECT 106.740 104.220 106.910 104.390 ;
        RECT 104.020 104.190 105.480 104.220 ;
        RECT 103.510 103.875 105.480 104.190 ;
        RECT 102.440 103.610 103.110 103.780 ;
        RECT 102.100 103.440 102.270 103.455 ;
        RECT 103.280 103.535 103.720 103.705 ;
        RECT 104.020 103.700 105.480 103.875 ;
        RECT 105.650 103.735 106.910 104.220 ;
        RECT 109.460 104.220 109.630 104.390 ;
        RECT 112.180 104.220 112.350 104.390 ;
        RECT 107.080 104.160 107.410 104.185 ;
        RECT 107.080 103.990 107.420 104.160 ;
        RECT 107.590 104.015 108.820 104.185 ;
        RECT 109.460 104.115 110.175 104.220 ;
        RECT 107.080 103.905 107.410 103.990 ;
        RECT 103.280 103.440 103.450 103.535 ;
        RECT 101.300 103.115 101.930 103.285 ;
        RECT 101.300 101.930 101.470 103.115 ;
        RECT 102.100 103.010 103.450 103.440 ;
        RECT 104.020 103.365 104.940 103.700 ;
        RECT 105.650 103.530 107.410 103.735 ;
        RECT 103.620 103.035 104.940 103.365 ;
        RECT 104.020 103.010 104.940 103.035 ;
        RECT 105.110 103.485 107.410 103.530 ;
        RECT 105.110 103.010 106.910 103.485 ;
        RECT 98.580 100.995 98.750 101.630 ;
        RECT 99.320 101.610 100.330 101.780 ;
        RECT 100.500 101.650 101.470 101.930 ;
        RECT 104.020 101.915 104.190 103.010 ;
        RECT 99.660 101.505 99.990 101.610 ;
        RECT 101.300 101.470 101.470 101.650 ;
        RECT 101.640 101.640 102.650 101.915 ;
        RECT 99.080 101.335 99.425 101.440 ;
        RECT 100.160 101.335 101.130 101.440 ;
        RECT 99.080 101.165 101.130 101.335 ;
        RECT 101.300 101.140 102.270 101.470 ;
        RECT 101.300 100.995 101.470 101.140 ;
        RECT 98.580 100.825 99.665 100.995 ;
        RECT 100.120 100.825 101.470 100.995 ;
        RECT 102.440 100.970 102.650 101.640 ;
        RECT 102.830 101.195 103.030 101.915 ;
        RECT 103.200 101.640 104.190 101.915 ;
        RECT 104.360 101.895 104.580 102.820 ;
        RECT 104.750 102.610 106.570 102.840 ;
        RECT 104.750 102.065 105.000 102.610 ;
        RECT 105.890 102.525 106.570 102.610 ;
        RECT 105.180 102.135 105.390 102.440 ;
        RECT 105.180 101.965 105.720 102.135 ;
        RECT 104.360 101.645 105.010 101.895 ;
        RECT 104.020 101.475 104.190 101.640 ;
        RECT 103.200 101.140 103.850 101.470 ;
        RECT 104.020 101.305 104.660 101.475 ;
        RECT 93.140 100.540 93.310 100.710 ;
        RECT 89.620 100.300 91.680 100.540 ;
        RECT 89.280 100.130 89.450 100.300 ;
        RECT 88.040 99.790 88.370 100.130 ;
        RECT 88.540 99.790 89.110 100.130 ;
        RECT 89.280 99.790 90.250 100.130 ;
        RECT 86.110 98.560 86.290 99.520 ;
        RECT 86.460 98.740 86.790 99.350 ;
        RECT 87.000 98.865 87.530 99.210 ;
        RECT 87.700 99.145 87.870 99.770 ;
        RECT 90.420 99.620 91.680 100.300 ;
        RECT 91.850 100.525 93.310 100.540 ;
        RECT 91.850 100.230 94.090 100.525 ;
        RECT 91.850 99.790 93.310 100.230 ;
        RECT 94.260 99.980 94.900 100.480 ;
        RECT 86.110 98.235 86.710 98.560 ;
        RECT 86.540 98.230 86.710 98.235 ;
        RECT 85.320 97.380 85.500 98.020 ;
        RECT 87.000 97.870 87.170 98.865 ;
        RECT 87.700 98.850 88.650 99.145 ;
        RECT 87.700 98.405 87.870 98.850 ;
        RECT 88.820 98.600 89.460 99.100 ;
        RECT 87.340 98.075 87.870 98.405 ;
        RECT 87.000 97.850 87.530 97.870 ;
        RECT 85.670 97.550 87.530 97.850 ;
        RECT 87.700 97.485 87.870 98.075 ;
        RECT 88.040 97.945 88.570 98.290 ;
        RECT 85.320 97.075 85.990 97.380 ;
        RECT 87.700 97.370 88.230 97.485 ;
        RECT 86.160 97.090 86.790 97.365 ;
        RECT 86.960 97.155 88.230 97.370 ;
        RECT 86.960 97.040 87.870 97.155 ;
        RECT 85.370 95.200 85.660 96.860 ;
        RECT 85.830 96.535 86.290 96.860 ;
        RECT 85.830 95.435 86.000 96.535 ;
        RECT 86.460 96.505 87.030 96.860 ;
        RECT 87.700 96.855 87.870 97.040 ;
        RECT 88.400 96.950 88.570 97.945 ;
        RECT 88.780 97.820 89.110 98.430 ;
        RECT 89.280 97.640 89.460 98.600 ;
        RECT 88.860 97.315 89.460 97.640 ;
        RECT 89.640 98.875 90.250 99.135 ;
        RECT 89.640 98.195 89.890 98.875 ;
        RECT 90.420 98.870 92.200 99.620 ;
        RECT 92.370 98.870 93.310 99.790 ;
        RECT 93.480 99.325 94.010 99.670 ;
        RECT 90.420 98.705 90.590 98.870 ;
        RECT 90.060 98.375 90.590 98.705 ;
        RECT 89.640 98.025 90.250 98.195 ;
        RECT 89.640 97.430 89.810 98.025 ;
        RECT 90.420 97.770 90.590 98.375 ;
        RECT 93.140 98.865 93.310 98.870 ;
        RECT 93.140 98.535 93.670 98.865 ;
        RECT 89.980 97.600 90.590 97.770 ;
        RECT 88.860 97.310 89.030 97.315 ;
        RECT 89.640 97.100 90.250 97.430 ;
        RECT 87.200 96.520 87.870 96.855 ;
        RECT 88.040 96.930 88.570 96.950 ;
        RECT 88.040 96.630 89.900 96.930 ;
        RECT 87.700 96.450 87.870 96.520 ;
        RECT 90.070 96.460 90.250 97.100 ;
        RECT 86.170 96.335 86.340 96.340 ;
        RECT 86.170 95.625 86.790 96.335 ;
        RECT 86.960 96.150 87.480 96.320 ;
        RECT 85.830 95.265 86.290 95.435 ;
        RECT 84.600 95.030 85.150 95.195 ;
        RECT 84.600 94.865 85.950 95.030 ;
        RECT 84.980 94.750 85.950 94.865 ;
        RECT 86.120 94.880 86.290 95.265 ;
        RECT 86.460 95.050 86.790 95.455 ;
        RECT 86.960 95.450 87.130 96.150 ;
        RECT 87.700 96.120 88.610 96.450 ;
        RECT 88.780 96.170 89.410 96.445 ;
        RECT 89.580 96.155 90.250 96.460 ;
        RECT 90.420 96.410 90.590 97.600 ;
        RECT 90.810 96.580 91.100 98.240 ;
        RECT 91.270 97.915 91.730 98.240 ;
        RECT 91.270 96.815 91.440 97.915 ;
        RECT 91.900 97.885 92.470 98.240 ;
        RECT 93.140 98.235 93.310 98.535 ;
        RECT 93.840 98.330 94.010 99.325 ;
        RECT 94.220 99.200 94.550 99.810 ;
        RECT 94.720 99.020 94.900 99.980 ;
        RECT 94.300 98.695 94.900 99.020 ;
        RECT 95.080 100.255 95.690 100.515 ;
        RECT 95.080 99.575 95.330 100.255 ;
        RECT 95.860 100.085 96.030 100.710 ;
        RECT 96.200 100.480 96.530 100.505 ;
        RECT 96.200 100.310 96.540 100.480 ;
        RECT 96.710 100.335 97.940 100.505 ;
        RECT 98.580 100.490 98.750 100.825 ;
        RECT 98.580 100.435 99.220 100.490 ;
        RECT 96.200 100.225 96.530 100.310 ;
        RECT 95.500 100.055 96.030 100.085 ;
        RECT 95.500 99.805 96.530 100.055 ;
        RECT 95.500 99.755 96.030 99.805 ;
        RECT 95.080 99.405 95.690 99.575 ;
        RECT 95.080 98.810 95.250 99.405 ;
        RECT 95.860 99.150 96.030 99.755 ;
        RECT 95.420 98.980 96.030 99.150 ;
        RECT 94.300 98.690 94.470 98.695 ;
        RECT 95.080 98.480 95.690 98.810 ;
        RECT 92.640 97.900 93.310 98.235 ;
        RECT 93.480 98.310 94.010 98.330 ;
        RECT 93.480 98.010 95.340 98.310 ;
        RECT 93.140 97.830 93.310 97.900 ;
        RECT 95.510 97.840 95.690 98.480 ;
        RECT 91.610 97.005 92.230 97.715 ;
        RECT 92.400 97.530 92.920 97.700 ;
        RECT 91.270 96.645 91.730 96.815 ;
        RECT 90.420 96.130 91.390 96.410 ;
        RECT 91.560 96.260 91.730 96.645 ;
        RECT 91.900 96.430 92.230 96.835 ;
        RECT 92.400 96.830 92.570 97.530 ;
        RECT 93.140 97.500 94.050 97.830 ;
        RECT 94.220 97.550 94.850 97.825 ;
        RECT 95.020 97.535 95.690 97.840 ;
        RECT 95.860 97.855 96.030 98.980 ;
        RECT 96.200 99.560 96.530 99.635 ;
        RECT 96.200 99.390 96.540 99.560 ;
        RECT 96.200 99.385 96.530 99.390 ;
        RECT 96.200 98.795 96.370 99.385 ;
        RECT 96.710 99.215 96.880 100.335 ;
        RECT 97.760 100.095 97.940 100.335 ;
        RECT 98.110 100.265 99.220 100.435 ;
        RECT 98.580 100.200 99.220 100.265 ;
        RECT 99.400 100.245 100.330 100.460 ;
        RECT 97.390 99.920 97.590 100.080 ;
        RECT 96.540 98.965 96.880 99.215 ;
        RECT 96.200 98.545 96.530 98.795 ;
        RECT 96.710 98.575 96.880 98.965 ;
        RECT 97.050 99.750 97.590 99.920 ;
        RECT 97.760 99.765 98.410 100.095 ;
        RECT 97.050 98.915 97.220 99.750 ;
        RECT 97.390 99.085 97.590 99.580 ;
        RECT 97.760 99.255 97.940 99.765 ;
        RECT 98.580 99.595 98.750 100.200 ;
        RECT 99.400 100.030 99.570 100.245 ;
        RECT 98.920 99.700 99.570 100.030 ;
        RECT 98.110 99.530 98.750 99.595 ;
        RECT 98.110 99.425 99.220 99.530 ;
        RECT 98.580 99.360 99.220 99.425 ;
        RECT 97.760 98.925 98.410 99.255 ;
        RECT 97.050 98.745 97.590 98.915 ;
        RECT 98.580 98.755 98.750 99.360 ;
        RECT 99.390 99.190 99.570 99.700 ;
        RECT 99.740 99.305 99.940 100.075 ;
        RECT 100.110 100.030 100.330 100.245 ;
        RECT 100.500 100.200 101.130 100.500 ;
        RECT 100.110 99.700 100.790 100.030 ;
        RECT 100.960 99.530 101.130 100.200 ;
        RECT 100.120 99.360 101.130 99.530 ;
        RECT 101.300 99.620 101.470 100.825 ;
        RECT 101.640 100.800 102.650 100.970 ;
        RECT 101.640 100.130 101.810 100.800 ;
        RECT 101.980 100.300 102.660 100.630 ;
        RECT 101.640 99.830 102.270 100.130 ;
        RECT 102.440 100.085 102.660 100.300 ;
        RECT 102.830 100.255 103.030 101.025 ;
        RECT 103.200 100.630 103.380 101.140 ;
        RECT 104.020 100.970 104.190 101.305 ;
        RECT 104.830 101.135 105.010 101.645 ;
        RECT 103.550 100.800 104.190 100.970 ;
        RECT 104.360 100.805 105.010 101.135 ;
        RECT 103.200 100.300 103.850 100.630 ;
        RECT 104.020 100.495 104.190 100.800 ;
        RECT 104.020 100.325 105.010 100.495 ;
        RECT 103.200 100.085 103.370 100.300 ;
        RECT 104.020 100.130 104.190 100.325 ;
        RECT 105.180 100.220 105.380 101.670 ;
        RECT 102.440 99.870 103.370 100.085 ;
        RECT 102.490 99.850 102.660 99.870 ;
        RECT 103.550 99.840 104.190 100.130 ;
        RECT 104.020 99.655 104.190 99.840 ;
        RECT 104.360 99.825 105.010 100.155 ;
        RECT 105.550 99.995 105.720 101.965 ;
        RECT 104.020 99.620 104.660 99.655 ;
        RECT 98.920 98.860 99.570 99.190 ;
        RECT 96.710 98.405 97.220 98.575 ;
        RECT 96.200 98.235 96.540 98.340 ;
        RECT 96.200 98.025 96.880 98.235 ;
        RECT 95.860 97.605 96.530 97.855 ;
        RECT 93.140 97.330 93.310 97.500 ;
        RECT 92.740 97.230 93.310 97.330 ;
        RECT 95.860 97.230 96.030 97.605 ;
        RECT 96.710 97.435 96.880 98.025 ;
        RECT 92.740 97.000 93.790 97.230 ;
        RECT 93.140 96.930 93.790 97.000 ;
        RECT 92.400 96.660 92.920 96.830 ;
        RECT 92.400 96.260 92.570 96.660 ;
        RECT 93.140 96.490 93.310 96.930 ;
        RECT 93.960 96.790 94.945 97.230 ;
        RECT 95.115 97.015 96.030 97.230 ;
        RECT 96.200 97.185 96.880 97.435 ;
        RECT 95.115 96.960 96.530 97.015 ;
        RECT 93.960 96.760 95.685 96.790 ;
        RECT 93.505 96.500 95.685 96.760 ;
        RECT 95.860 96.710 96.530 96.960 ;
        RECT 87.700 95.950 87.870 96.120 ;
        RECT 87.300 95.935 87.870 95.950 ;
        RECT 87.300 95.620 88.370 95.935 ;
        RECT 87.700 95.600 88.370 95.620 ;
        RECT 86.960 95.280 87.480 95.450 ;
        RECT 86.960 94.880 87.130 95.280 ;
        RECT 87.700 95.110 87.870 95.600 ;
        RECT 88.540 95.585 89.110 95.940 ;
        RECT 89.280 95.615 89.740 95.940 ;
        RECT 89.230 95.415 89.400 95.420 ;
        RECT 88.090 95.230 88.610 95.400 ;
        RECT 84.260 94.270 84.810 94.695 ;
        RECT 80.390 93.980 80.580 94.120 ;
        RECT 79.105 93.790 80.580 93.980 ;
        RECT 80.750 93.905 82.040 94.160 ;
        RECT 79.105 93.355 80.215 93.790 ;
        RECT 80.750 93.620 80.920 93.905 ;
        RECT 80.385 93.365 80.920 93.620 ;
        RECT 76.275 92.435 76.990 93.355 ;
        RECT 74.095 92.360 74.270 92.435 ;
        RECT 73.370 92.115 74.270 92.360 ;
        RECT 72.960 91.685 73.925 91.945 ;
        RECT 74.095 91.800 74.270 92.115 ;
        RECT 76.820 91.800 76.990 92.435 ;
        RECT 79.540 93.350 80.215 93.355 ;
        RECT 81.100 93.350 81.580 93.735 ;
        RECT 81.775 93.370 82.040 93.905 ;
        RECT 79.540 93.180 79.710 93.350 ;
        RECT 82.260 93.180 82.430 94.270 ;
        RECT 84.980 94.095 85.150 94.750 ;
        RECT 86.120 94.710 87.130 94.880 ;
        RECT 87.300 95.030 87.870 95.110 ;
        RECT 87.300 94.730 88.270 95.030 ;
        RECT 86.460 94.605 86.790 94.710 ;
        RECT 87.700 94.700 88.270 94.730 ;
        RECT 85.320 94.435 86.290 94.540 ;
        RECT 87.025 94.435 87.370 94.540 ;
        RECT 85.320 94.265 87.370 94.435 ;
        RECT 87.700 94.190 87.870 94.700 ;
        RECT 88.440 94.530 88.610 95.230 ;
        RECT 88.780 94.705 89.400 95.415 ;
        RECT 88.090 94.360 88.610 94.530 ;
        RECT 87.700 94.095 88.270 94.190 ;
        RECT 84.980 93.925 86.330 94.095 ;
        RECT 86.785 93.925 88.270 94.095 ;
        RECT 84.980 93.640 85.150 93.925 ;
        RECT 87.700 93.810 88.270 93.925 ;
        RECT 88.440 93.960 88.610 94.360 ;
        RECT 88.780 94.130 89.110 94.535 ;
        RECT 89.570 94.515 89.740 95.615 ;
        RECT 89.280 94.345 89.740 94.515 ;
        RECT 89.280 93.960 89.450 94.345 ;
        RECT 89.910 94.280 90.200 95.940 ;
        RECT 90.420 95.475 90.590 96.130 ;
        RECT 91.560 96.090 92.570 96.260 ;
        RECT 92.740 96.330 93.310 96.490 ;
        RECT 92.740 96.110 93.790 96.330 ;
        RECT 91.900 95.985 92.230 96.090 ;
        RECT 93.140 96.070 93.790 96.110 ;
        RECT 90.760 95.815 91.730 95.920 ;
        RECT 92.465 95.815 92.810 95.920 ;
        RECT 90.760 95.645 92.810 95.815 ;
        RECT 93.140 95.475 93.310 96.070 ;
        RECT 93.960 96.065 94.945 96.500 ;
        RECT 95.860 96.330 96.030 96.710 ;
        RECT 96.710 96.540 96.880 97.185 ;
        RECT 95.130 96.075 96.030 96.330 ;
        RECT 93.960 95.890 94.130 96.065 ;
        RECT 93.505 95.630 94.130 95.890 ;
        RECT 90.420 95.305 91.770 95.475 ;
        RECT 92.225 95.460 93.310 95.475 ;
        RECT 92.225 95.305 93.790 95.460 ;
        RECT 90.420 94.110 90.590 95.305 ;
        RECT 93.140 95.210 93.790 95.305 ;
        RECT 87.700 93.640 87.870 93.810 ;
        RECT 88.440 93.790 89.450 93.960 ;
        RECT 89.620 93.830 90.590 94.110 ;
        RECT 88.780 93.685 89.110 93.790 ;
        RECT 79.540 92.490 80.800 93.180 ;
        RECT 80.970 92.660 82.430 93.180 ;
        RECT 72.960 91.085 73.200 91.685 ;
        RECT 74.095 91.515 75.435 91.800 ;
        RECT 73.370 91.510 75.435 91.515 ;
        RECT 76.095 91.510 76.990 91.800 ;
        RECT 73.370 91.340 74.270 91.510 ;
        RECT 76.820 91.340 76.990 91.510 ;
        RECT 73.370 91.255 75.280 91.340 ;
        RECT 72.960 90.825 73.925 91.085 ;
        RECT 74.095 91.080 75.280 91.255 ;
        RECT 72.960 90.225 73.200 90.825 ;
        RECT 74.095 90.655 74.270 91.080 ;
        RECT 75.460 90.910 75.980 91.340 ;
        RECT 76.160 91.065 76.990 91.340 ;
        RECT 77.160 91.315 77.380 92.240 ;
        RECT 77.550 92.030 79.370 92.260 ;
        RECT 77.550 91.485 77.800 92.030 ;
        RECT 78.690 91.945 79.370 92.030 ;
        RECT 79.540 91.970 81.340 92.490 ;
        RECT 81.510 91.970 82.430 92.660 ;
        RECT 82.600 92.235 82.820 93.160 ;
        RECT 82.990 92.950 84.810 93.180 ;
        RECT 82.990 92.405 83.240 92.950 ;
        RECT 84.130 92.865 84.810 92.950 ;
        RECT 83.420 92.475 83.630 92.780 ;
        RECT 83.420 92.305 83.960 92.475 ;
        RECT 82.600 91.985 83.250 92.235 ;
        RECT 77.980 91.555 78.190 91.860 ;
        RECT 77.980 91.385 78.520 91.555 ;
        RECT 77.160 91.065 77.810 91.315 ;
        RECT 73.370 90.435 74.270 90.655 ;
        RECT 74.440 90.895 75.980 90.910 ;
        RECT 76.820 90.895 76.990 91.065 ;
        RECT 74.440 90.740 76.650 90.895 ;
        RECT 74.440 90.635 75.110 90.740 ;
        RECT 75.460 90.725 76.650 90.740 ;
        RECT 76.190 90.645 76.650 90.725 ;
        RECT 76.820 90.725 77.460 90.895 ;
        RECT 73.370 90.395 75.115 90.435 ;
        RECT 72.960 89.965 73.925 90.225 ;
        RECT 74.095 90.220 75.115 90.395 ;
        RECT 75.310 90.325 75.910 90.555 ;
        RECT 76.820 90.470 76.990 90.725 ;
        RECT 77.630 90.555 77.810 91.065 ;
        RECT 72.960 89.365 73.200 89.965 ;
        RECT 74.095 89.795 74.270 90.220 ;
        RECT 73.370 89.535 74.270 89.795 ;
        RECT 74.440 89.560 74.780 90.035 ;
        RECT 75.310 89.995 75.480 90.325 ;
        RECT 76.325 90.140 76.990 90.470 ;
        RECT 77.160 90.225 77.810 90.555 ;
        RECT 75.015 89.745 75.480 89.995 ;
        RECT 75.310 89.560 75.480 89.745 ;
        RECT 75.660 89.960 76.155 90.140 ;
        RECT 75.660 89.730 76.600 89.960 ;
        RECT 76.820 89.915 76.990 90.140 ;
        RECT 76.820 89.745 77.810 89.915 ;
        RECT 74.095 89.380 74.270 89.535 ;
        RECT 74.950 89.380 75.140 89.520 ;
        RECT 72.960 89.105 73.925 89.365 ;
        RECT 74.095 89.190 75.140 89.380 ;
        RECT 75.310 89.305 76.600 89.560 ;
        RECT 74.095 88.935 74.775 89.190 ;
        RECT 75.310 89.020 75.480 89.305 ;
        RECT 73.300 88.750 74.775 88.935 ;
        RECT 74.945 88.765 75.480 89.020 ;
        RECT 75.660 88.750 76.140 89.135 ;
        RECT 76.335 88.770 76.600 89.305 ;
        RECT 76.820 89.075 76.990 89.745 ;
        RECT 77.980 89.640 78.180 91.090 ;
        RECT 77.160 89.245 77.810 89.575 ;
        RECT 78.350 89.415 78.520 91.385 ;
        RECT 76.820 88.905 77.460 89.075 ;
        RECT 73.300 88.675 74.270 88.750 ;
        RECT 74.100 88.580 74.270 88.675 ;
        RECT 76.820 88.580 76.990 88.905 ;
        RECT 77.630 88.735 77.810 89.245 ;
        RECT 62.785 87.880 63.850 88.145 ;
        RECT 64.360 87.935 65.310 88.215 ;
        RECT 65.940 88.130 66.110 88.250 ;
        RECT 65.480 87.880 66.110 88.130 ;
        RECT 60.500 87.115 62.045 87.455 ;
        RECT 60.500 83.695 61.215 87.115 ;
        RECT 62.785 85.975 63.390 87.880 ;
        RECT 63.985 87.710 65.350 87.765 ;
        RECT 63.560 87.595 65.660 87.710 ;
        RECT 63.560 87.460 64.115 87.595 ;
        RECT 65.220 87.540 65.660 87.595 ;
        RECT 63.665 86.315 63.835 87.250 ;
        RECT 64.305 87.185 64.900 87.425 ;
        RECT 65.490 87.375 65.660 87.540 ;
        RECT 65.070 87.015 65.290 87.370 ;
        RECT 64.005 86.845 65.290 87.015 ;
        RECT 64.005 86.485 64.370 86.845 ;
        RECT 65.490 86.675 65.660 87.180 ;
        RECT 64.540 86.505 65.660 86.675 ;
        RECT 65.940 86.900 66.110 87.880 ;
        RECT 66.390 87.685 67.350 88.065 ;
        RECT 67.695 87.630 67.960 88.300 ;
        RECT 68.660 88.130 68.830 88.340 ;
        RECT 69.425 88.170 70.790 88.225 ;
        RECT 68.150 87.800 68.830 88.130 ;
        RECT 69.000 88.055 71.100 88.170 ;
        RECT 69.000 87.920 69.555 88.055 ;
        RECT 70.660 88.000 71.100 88.055 ;
        RECT 67.695 87.405 68.490 87.630 ;
        RECT 66.280 87.120 66.850 87.310 ;
        RECT 65.940 86.570 66.470 86.900 ;
        RECT 66.680 86.740 66.850 87.120 ;
        RECT 67.020 86.910 67.435 87.235 ;
        RECT 67.715 86.920 68.490 87.235 ;
        RECT 67.715 86.740 67.945 86.920 ;
        RECT 66.680 86.570 67.945 86.740 ;
        RECT 68.660 86.730 68.830 87.800 ;
        RECT 64.540 86.315 64.710 86.505 ;
        RECT 63.665 86.145 64.710 86.315 ;
        RECT 64.450 85.975 64.710 86.145 ;
        RECT 64.930 86.095 65.260 86.295 ;
        RECT 65.940 86.185 66.110 86.570 ;
        RECT 67.020 86.400 67.945 86.570 ;
        RECT 68.245 86.435 68.830 86.730 ;
        RECT 69.105 86.775 69.275 87.710 ;
        RECT 69.745 87.645 70.340 87.885 ;
        RECT 70.930 87.835 71.100 88.000 ;
        RECT 71.380 88.075 71.550 88.340 ;
        RECT 71.730 88.255 73.925 88.505 ;
        RECT 70.510 87.475 70.730 87.830 ;
        RECT 71.380 87.815 72.075 88.075 ;
        RECT 69.445 87.305 70.730 87.475 ;
        RECT 69.445 86.945 69.810 87.305 ;
        RECT 70.930 87.135 71.100 87.640 ;
        RECT 69.980 86.965 71.100 87.135 ;
        RECT 71.380 87.215 71.550 87.815 ;
        RECT 72.540 87.645 72.790 88.255 ;
        RECT 74.100 88.075 74.705 88.580 ;
        RECT 73.290 87.815 74.705 88.075 ;
        RECT 71.730 87.640 72.790 87.645 ;
        RECT 71.730 87.395 73.930 87.640 ;
        RECT 69.980 86.775 70.150 86.965 ;
        RECT 69.105 86.605 70.150 86.775 ;
        RECT 71.380 86.910 72.060 87.215 ;
        RECT 72.230 86.910 72.790 87.225 ;
        RECT 74.100 87.215 74.705 87.815 ;
        RECT 73.290 86.920 74.705 87.215 ;
        RECT 76.275 88.200 76.990 88.580 ;
        RECT 77.160 88.370 77.810 88.735 ;
        RECT 77.980 89.245 78.520 89.415 ;
        RECT 78.690 91.355 78.870 91.945 ;
        RECT 79.540 91.800 79.710 91.970 ;
        RECT 82.260 91.815 82.430 91.970 ;
        RECT 82.260 91.800 82.900 91.815 ;
        RECT 79.540 91.775 80.875 91.800 ;
        RECT 79.040 91.525 80.875 91.775 ;
        RECT 79.540 91.510 80.875 91.525 ;
        RECT 81.535 91.645 82.900 91.800 ;
        RECT 81.535 91.510 82.430 91.645 ;
        RECT 78.690 91.105 79.370 91.355 ;
        RECT 79.540 91.160 79.710 91.510 ;
        RECT 82.260 91.170 82.430 91.510 ;
        RECT 83.070 91.475 83.250 91.985 ;
        RECT 78.690 90.515 78.870 91.105 ;
        RECT 79.540 90.990 80.625 91.160 ;
        RECT 81.745 91.000 82.430 91.170 ;
        RECT 82.600 91.145 83.250 91.475 ;
        RECT 79.540 90.935 79.710 90.990 ;
        RECT 79.040 90.685 79.710 90.935 ;
        RECT 80.770 90.830 81.605 90.880 ;
        RECT 82.260 90.835 82.430 91.000 ;
        RECT 80.770 90.820 82.040 90.830 ;
        RECT 78.690 90.265 79.370 90.515 ;
        RECT 79.540 90.320 79.710 90.685 ;
        RECT 79.925 90.710 82.040 90.820 ;
        RECT 79.925 90.665 80.900 90.710 ;
        RECT 79.925 90.490 80.850 90.665 ;
        RECT 81.480 90.655 82.040 90.710 ;
        RECT 77.980 88.390 78.190 89.245 ;
        RECT 78.690 89.035 78.860 90.265 ;
        RECT 79.540 90.150 80.720 90.320 ;
        RECT 79.030 89.705 79.370 89.955 ;
        RECT 79.540 89.535 79.710 90.150 ;
        RECT 81.020 89.990 81.350 90.540 ;
        RECT 81.520 90.500 82.040 90.655 ;
        RECT 82.260 90.665 83.250 90.835 ;
        RECT 82.260 90.330 82.430 90.665 ;
        RECT 83.420 90.560 83.620 92.010 ;
        RECT 81.650 90.160 82.430 90.330 ;
        RECT 82.600 90.165 83.250 90.495 ;
        RECT 83.790 90.335 83.960 92.305 ;
        RECT 82.260 89.995 82.430 90.160 ;
        RECT 81.020 89.980 82.045 89.990 ;
        RECT 79.880 89.790 82.045 89.980 ;
        RECT 79.880 89.640 80.815 89.790 ;
        RECT 81.520 89.660 82.045 89.790 ;
        RECT 82.260 89.825 82.900 89.995 ;
        RECT 79.040 89.410 79.710 89.535 ;
        RECT 79.040 89.285 80.210 89.410 ;
        RECT 78.360 88.865 78.860 89.035 ;
        RECT 76.275 88.030 77.460 88.200 ;
        RECT 76.275 86.995 76.990 88.030 ;
        RECT 69.890 86.435 70.150 86.605 ;
        RECT 70.370 86.555 70.700 86.755 ;
        RECT 71.380 86.740 71.550 86.910 ;
        RECT 74.100 86.740 74.705 86.920 ;
        RECT 71.380 86.645 72.210 86.740 ;
        RECT 68.245 86.400 69.630 86.435 ;
        RECT 66.280 86.230 66.850 86.400 ;
        RECT 68.660 86.265 69.630 86.400 ;
        RECT 69.890 86.265 70.220 86.435 ;
        RECT 66.280 86.210 68.490 86.230 ;
        RECT 62.785 85.805 64.190 85.975 ;
        RECT 64.450 85.805 64.780 85.975 ;
        RECT 62.785 85.635 63.390 85.805 ;
        RECT 64.960 85.635 65.260 86.095 ;
        RECT 65.440 86.040 66.110 86.185 ;
        RECT 65.440 85.815 66.490 86.040 ;
        RECT 66.660 86.000 68.490 86.210 ;
        RECT 68.660 85.830 68.830 86.265 ;
        RECT 70.400 86.095 70.700 86.555 ;
        RECT 70.880 86.465 72.210 86.645 ;
        RECT 70.880 86.275 71.550 86.465 ;
        RECT 72.390 86.310 72.910 86.740 ;
        RECT 73.090 86.480 74.705 86.740 ;
        RECT 75.445 86.655 76.990 86.995 ;
        RECT 72.390 86.295 73.930 86.310 ;
        RECT 69.000 85.925 71.100 86.095 ;
        RECT 69.000 85.845 69.330 85.925 ;
        RECT 65.940 85.710 66.490 85.815 ;
        RECT 61.535 85.285 63.390 85.635 ;
        RECT 63.560 85.465 65.660 85.635 ;
        RECT 63.560 85.385 63.890 85.465 ;
        RECT 62.785 84.095 63.390 85.285 ;
        RECT 63.690 84.445 63.860 85.160 ;
        RECT 64.060 85.105 64.780 85.295 ;
        RECT 65.490 85.230 65.660 85.465 ;
        RECT 65.940 85.360 66.110 85.710 ;
        RECT 67.690 85.540 68.830 85.830 ;
        RECT 68.660 85.360 68.830 85.540 ;
        RECT 64.990 84.935 65.320 85.080 ;
        RECT 64.030 84.615 65.320 84.935 ;
        RECT 65.490 84.445 65.660 85.060 ;
        RECT 63.690 84.275 65.660 84.445 ;
        RECT 65.940 84.840 67.400 85.360 ;
        RECT 62.785 83.780 63.890 84.095 ;
        RECT 62.785 83.695 63.390 83.780 ;
        RECT 60.500 83.520 60.670 83.695 ;
        RECT 63.220 83.520 63.390 83.695 ;
        RECT 64.120 83.550 64.495 84.105 ;
        RECT 64.700 83.570 65.030 84.275 ;
        RECT 65.940 84.150 66.860 84.840 ;
        RECT 67.570 84.670 68.830 85.360 ;
        RECT 69.130 84.905 69.300 85.620 ;
        RECT 69.500 85.565 70.220 85.755 ;
        RECT 70.930 85.690 71.100 85.925 ;
        RECT 71.380 85.870 71.550 86.275 ;
        RECT 71.720 86.140 73.930 86.295 ;
        RECT 71.720 86.125 72.910 86.140 ;
        RECT 71.720 86.045 72.180 86.125 ;
        RECT 73.260 86.035 73.930 86.140 ;
        RECT 71.380 85.540 72.045 85.870 ;
        RECT 72.460 85.725 73.060 85.955 ;
        RECT 74.100 85.835 74.705 86.480 ;
        RECT 70.430 85.395 70.760 85.540 ;
        RECT 69.470 85.075 70.760 85.395 ;
        RECT 70.930 84.905 71.100 85.520 ;
        RECT 69.130 84.735 71.100 84.905 ;
        RECT 67.030 84.555 68.830 84.670 ;
        RECT 67.030 84.240 69.330 84.555 ;
        RECT 67.030 84.150 68.830 84.240 ;
        RECT 65.940 84.000 66.110 84.150 ;
        RECT 65.410 83.790 66.110 84.000 ;
        RECT 68.660 83.970 68.830 84.150 ;
        RECT 69.560 84.010 69.935 84.565 ;
        RECT 70.140 84.030 70.470 84.735 ;
        RECT 71.380 84.460 71.550 85.540 ;
        RECT 72.215 85.360 72.710 85.540 ;
        RECT 71.770 85.130 72.710 85.360 ;
        RECT 72.890 85.395 73.060 85.725 ;
        RECT 73.255 85.620 74.705 85.835 ;
        RECT 72.890 85.145 73.355 85.395 ;
        RECT 72.890 84.960 73.060 85.145 ;
        RECT 73.590 84.960 73.930 85.435 ;
        RECT 74.100 85.175 74.705 85.620 ;
        RECT 76.275 86.280 76.990 86.655 ;
        RECT 77.210 86.840 77.380 87.760 ;
        RECT 77.630 87.340 77.810 88.370 ;
        RECT 78.360 87.710 78.530 88.865 ;
        RECT 79.030 88.790 79.370 89.115 ;
        RECT 77.550 87.010 77.810 87.340 ;
        RECT 77.980 87.540 78.530 87.710 ;
        RECT 78.700 88.410 79.030 88.620 ;
        RECT 77.980 87.050 78.150 87.540 ;
        RECT 78.700 87.300 78.870 88.410 ;
        RECT 79.200 88.240 79.370 88.790 ;
        RECT 79.040 87.990 79.370 88.240 ;
        RECT 79.540 89.095 80.210 89.285 ;
        RECT 79.540 87.720 79.710 89.095 ;
        RECT 80.440 89.085 80.815 89.640 ;
        RECT 81.020 88.915 81.350 89.620 ;
        RECT 82.260 89.400 82.430 89.825 ;
        RECT 83.070 89.655 83.250 90.165 ;
        RECT 81.730 89.190 82.430 89.400 ;
        RECT 82.600 89.290 83.250 89.655 ;
        RECT 83.420 90.165 83.960 90.335 ;
        RECT 84.130 92.275 84.310 92.865 ;
        RECT 84.980 92.720 86.240 93.640 ;
        RECT 86.410 93.175 87.870 93.640 ;
        RECT 88.200 93.515 88.545 93.620 ;
        RECT 89.280 93.515 90.250 93.620 ;
        RECT 88.200 93.345 90.250 93.515 ;
        RECT 90.420 93.190 90.590 93.830 ;
        RECT 90.810 93.360 91.100 95.020 ;
        RECT 91.270 94.695 91.730 95.020 ;
        RECT 91.270 93.595 91.440 94.695 ;
        RECT 91.900 94.665 92.470 95.020 ;
        RECT 93.140 95.015 93.310 95.210 ;
        RECT 93.960 95.030 94.130 95.630 ;
        RECT 92.640 94.680 93.310 95.015 ;
        RECT 93.505 94.770 94.130 95.030 ;
        RECT 93.140 94.600 93.310 94.680 ;
        RECT 91.610 93.785 92.230 94.495 ;
        RECT 92.400 94.310 92.920 94.480 ;
        RECT 93.140 94.350 93.790 94.600 ;
        RECT 91.270 93.425 91.730 93.595 ;
        RECT 90.420 93.175 91.390 93.190 ;
        RECT 86.410 93.005 88.785 93.175 ;
        RECT 89.240 93.005 91.390 93.175 ;
        RECT 86.410 92.890 87.870 93.005 ;
        RECT 86.930 92.720 87.870 92.890 ;
        RECT 90.420 92.910 91.390 93.005 ;
        RECT 91.560 93.040 91.730 93.425 ;
        RECT 91.900 93.210 92.230 93.615 ;
        RECT 92.400 93.610 92.570 94.310 ;
        RECT 93.140 94.110 93.310 94.350 ;
        RECT 93.960 94.170 94.130 94.770 ;
        RECT 92.740 93.780 93.310 94.110 ;
        RECT 93.505 93.910 94.130 94.170 ;
        RECT 93.140 93.740 93.310 93.780 ;
        RECT 92.400 93.440 92.920 93.610 ;
        RECT 93.140 93.495 93.790 93.740 ;
        RECT 92.400 93.040 92.570 93.440 ;
        RECT 93.140 93.270 93.310 93.495 ;
        RECT 93.960 93.325 94.130 93.910 ;
        RECT 90.420 92.720 90.590 92.910 ;
        RECT 91.560 92.870 92.570 93.040 ;
        RECT 92.740 92.890 93.310 93.270 ;
        RECT 93.505 93.050 94.130 93.325 ;
        RECT 93.140 92.880 93.310 92.890 ;
        RECT 91.900 92.765 92.230 92.870 ;
        RECT 84.980 92.695 86.760 92.720 ;
        RECT 84.480 92.445 86.760 92.695 ;
        RECT 84.130 92.025 84.810 92.275 ;
        RECT 84.130 91.435 84.310 92.025 ;
        RECT 84.980 91.970 86.760 92.445 ;
        RECT 86.930 92.200 89.160 92.720 ;
        RECT 89.330 92.255 90.590 92.720 ;
        RECT 90.760 92.595 91.730 92.700 ;
        RECT 92.465 92.595 92.810 92.700 ;
        RECT 90.760 92.425 92.810 92.595 ;
        RECT 93.140 92.635 93.790 92.880 ;
        RECT 93.140 92.255 93.310 92.635 ;
        RECT 93.960 92.465 94.130 93.050 ;
        RECT 86.930 91.970 88.620 92.200 ;
        RECT 89.330 92.085 91.770 92.255 ;
        RECT 92.225 92.085 93.310 92.255 ;
        RECT 93.505 92.205 94.130 92.465 ;
        RECT 89.330 92.030 90.590 92.085 ;
        RECT 84.980 91.855 85.150 91.970 ;
        RECT 84.480 91.800 85.150 91.855 ;
        RECT 87.700 91.800 88.620 91.970 ;
        RECT 84.480 91.605 86.315 91.800 ;
        RECT 84.980 91.510 86.315 91.605 ;
        RECT 86.975 91.510 88.620 91.800 ;
        RECT 88.790 91.800 90.590 92.030 ;
        RECT 93.140 92.035 93.310 92.085 ;
        RECT 93.140 91.800 93.790 92.035 ;
        RECT 88.790 91.510 91.755 91.800 ;
        RECT 92.415 91.775 93.790 91.800 ;
        RECT 92.415 91.510 93.310 91.775 ;
        RECT 93.960 91.605 94.130 92.205 ;
        RECT 84.130 91.185 84.810 91.435 ;
        RECT 84.980 91.330 85.150 91.510 ;
        RECT 87.700 91.340 87.870 91.510 ;
        RECT 90.420 91.340 90.590 91.510 ;
        RECT 83.420 89.310 83.630 90.165 ;
        RECT 84.130 89.955 84.300 91.185 ;
        RECT 84.980 91.035 85.960 91.330 ;
        RECT 84.470 90.625 84.810 90.875 ;
        RECT 84.980 90.455 85.150 91.035 ;
        RECT 86.460 91.025 87.020 91.340 ;
        RECT 87.190 91.335 87.870 91.340 ;
        RECT 87.190 91.035 88.370 91.335 ;
        RECT 87.700 91.000 88.370 91.035 ;
        RECT 85.320 90.610 87.520 90.855 ;
        RECT 84.480 90.435 85.150 90.455 ;
        RECT 86.460 90.605 87.520 90.610 ;
        RECT 84.480 90.205 85.960 90.435 ;
        RECT 84.980 90.175 85.960 90.205 ;
        RECT 83.800 89.785 84.300 89.955 ;
        RECT 82.260 89.120 82.430 89.190 ;
        RECT 82.260 88.950 82.900 89.120 ;
        RECT 80.010 88.745 81.980 88.915 ;
        RECT 80.010 88.030 80.180 88.745 ;
        RECT 80.350 88.255 81.640 88.575 ;
        RECT 81.310 88.110 81.640 88.255 ;
        RECT 81.810 88.130 81.980 88.745 ;
        RECT 80.380 87.895 81.100 88.085 ;
        RECT 79.040 87.470 79.710 87.720 ;
        RECT 79.880 87.725 80.210 87.805 ;
        RECT 81.810 87.725 81.980 87.960 ;
        RECT 79.880 87.555 81.980 87.725 ;
        RECT 79.540 87.385 79.710 87.470 ;
        RECT 78.320 87.050 79.030 87.300 ;
        RECT 79.540 87.215 80.510 87.385 ;
        RECT 80.770 87.215 81.100 87.385 ;
        RECT 78.320 86.840 78.530 87.050 ;
        RECT 79.540 86.880 79.710 87.215 ;
        RECT 80.770 87.045 81.030 87.215 ;
        RECT 81.280 87.095 81.580 87.555 ;
        RECT 82.260 87.375 82.430 88.950 ;
        RECT 77.210 86.450 78.530 86.840 ;
        RECT 78.700 86.450 79.710 86.880 ;
        RECT 79.540 86.280 79.710 86.450 ;
        RECT 70.850 84.250 71.550 84.460 ;
        RECT 60.500 83.000 61.960 83.520 ;
        RECT 62.130 83.040 63.390 83.520 ;
        RECT 63.560 83.400 64.495 83.550 ;
        RECT 65.200 83.400 65.725 83.530 ;
        RECT 63.560 83.210 65.725 83.400 ;
        RECT 64.700 83.200 65.725 83.210 ;
        RECT 60.500 82.310 61.420 83.000 ;
        RECT 62.130 82.870 64.400 83.040 ;
        RECT 62.130 82.830 63.390 82.870 ;
        RECT 61.590 82.310 63.390 82.830 ;
        RECT 63.605 82.525 64.530 82.700 ;
        RECT 64.700 82.650 65.030 83.200 ;
        RECT 65.940 83.030 66.110 83.790 ;
        RECT 66.280 83.565 66.610 83.890 ;
        RECT 66.780 83.735 68.100 83.940 ;
        RECT 68.280 83.640 68.830 83.970 ;
        RECT 69.000 83.860 69.935 84.010 ;
        RECT 70.640 83.860 71.165 83.990 ;
        RECT 69.000 83.670 71.165 83.860 ;
        RECT 66.280 83.465 67.690 83.565 ;
        RECT 68.660 83.500 68.830 83.640 ;
        RECT 70.140 83.660 71.165 83.670 ;
        RECT 66.280 83.395 68.490 83.465 ;
        RECT 67.520 83.215 68.490 83.395 ;
        RECT 68.660 83.330 69.840 83.500 ;
        RECT 65.330 82.860 66.110 83.030 ;
        RECT 65.200 82.535 65.720 82.690 ;
        RECT 63.605 82.480 64.580 82.525 ;
        RECT 65.160 82.480 65.720 82.535 ;
        RECT 63.605 82.370 65.720 82.480 ;
        RECT 64.450 82.360 65.720 82.370 ;
        RECT 64.450 82.310 65.285 82.360 ;
        RECT 60.500 82.130 60.670 82.310 ;
        RECT 63.220 82.200 63.390 82.310 ;
        RECT 60.500 81.800 61.175 82.130 ;
        RECT 62.030 82.075 62.200 82.080 ;
        RECT 60.500 80.350 60.670 81.800 ;
        RECT 61.350 81.775 62.200 82.075 ;
        RECT 62.370 81.880 63.030 82.050 ;
        RECT 63.220 82.030 64.305 82.200 ;
        RECT 65.940 82.190 66.110 82.860 ;
        RECT 66.445 82.820 67.350 83.175 ;
        RECT 66.440 82.475 67.350 82.645 ;
        RECT 67.520 82.480 67.690 83.215 ;
        RECT 68.660 82.995 68.830 83.330 ;
        RECT 67.940 82.665 68.830 82.995 ;
        RECT 69.045 82.985 69.970 83.160 ;
        RECT 70.140 83.110 70.470 83.660 ;
        RECT 71.380 83.520 71.550 84.250 ;
        RECT 71.770 84.705 73.060 84.960 ;
        RECT 71.770 84.170 72.035 84.705 ;
        RECT 72.230 84.150 72.710 84.535 ;
        RECT 72.890 84.420 73.060 84.705 ;
        RECT 73.230 84.780 73.420 84.920 ;
        RECT 74.100 84.825 75.955 85.175 ;
        RECT 74.100 84.780 74.705 84.825 ;
        RECT 73.230 84.590 74.705 84.780 ;
        RECT 72.890 84.165 73.425 84.420 ;
        RECT 73.595 84.150 74.705 84.590 ;
        RECT 71.380 83.490 72.030 83.520 ;
        RECT 70.770 83.320 72.030 83.490 ;
        RECT 71.380 83.260 72.030 83.320 ;
        RECT 72.220 83.280 72.790 83.475 ;
        RECT 72.960 83.260 73.930 83.430 ;
        RECT 70.640 82.995 71.160 83.150 ;
        RECT 69.045 82.940 70.020 82.985 ;
        RECT 70.600 82.940 71.160 82.995 ;
        RECT 69.045 82.830 71.160 82.940 ;
        RECT 69.890 82.820 71.160 82.830 ;
        RECT 69.890 82.770 70.725 82.820 ;
        RECT 68.660 82.660 68.830 82.665 ;
        RECT 68.660 82.490 69.745 82.660 ;
        RECT 71.380 82.650 71.550 83.260 ;
        RECT 72.960 83.090 73.130 83.260 ;
        RECT 71.720 82.920 73.130 83.090 ;
        RECT 74.100 83.235 74.705 84.150 ;
        RECT 76.275 84.630 78.280 86.280 ;
        RECT 78.450 85.310 79.710 86.280 ;
        RECT 79.985 86.875 81.030 87.045 ;
        RECT 81.250 86.895 81.580 87.095 ;
        RECT 81.760 87.200 82.430 87.375 ;
        RECT 82.650 87.760 82.820 88.680 ;
        RECT 83.070 88.260 83.250 89.290 ;
        RECT 83.800 88.630 83.970 89.785 ;
        RECT 84.470 89.710 84.810 90.035 ;
        RECT 82.990 87.930 83.250 88.260 ;
        RECT 83.420 88.460 83.970 88.630 ;
        RECT 84.140 89.330 84.470 89.540 ;
        RECT 83.420 87.970 83.590 88.460 ;
        RECT 84.140 88.220 84.310 89.330 ;
        RECT 84.640 89.160 84.810 89.710 ;
        RECT 84.480 88.910 84.810 89.160 ;
        RECT 84.980 89.575 85.150 90.175 ;
        RECT 86.460 89.995 86.710 90.605 ;
        RECT 87.700 90.435 87.870 91.000 ;
        RECT 88.540 90.985 89.110 91.340 ;
        RECT 89.280 91.015 89.740 91.340 ;
        RECT 88.090 90.630 88.610 90.800 ;
        RECT 87.175 90.430 87.870 90.435 ;
        RECT 87.175 90.175 88.270 90.430 ;
        RECT 87.700 90.100 88.270 90.175 ;
        RECT 85.325 89.745 87.520 89.995 ;
        RECT 84.980 89.315 85.950 89.575 ;
        RECT 84.980 88.715 85.155 89.315 ;
        RECT 85.325 88.885 86.290 89.145 ;
        RECT 84.980 88.640 85.880 88.715 ;
        RECT 84.480 88.455 85.880 88.640 ;
        RECT 84.480 88.390 85.155 88.455 ;
        RECT 83.760 87.970 84.470 88.220 ;
        RECT 83.760 87.760 83.970 87.970 ;
        RECT 84.980 87.855 85.155 88.390 ;
        RECT 86.050 88.285 86.290 88.885 ;
        RECT 85.325 88.025 86.290 88.285 ;
        RECT 84.980 87.800 85.880 87.855 ;
        RECT 82.650 87.370 83.970 87.760 ;
        RECT 84.140 87.595 85.880 87.800 ;
        RECT 84.140 87.370 85.155 87.595 ;
        RECT 86.050 87.425 86.290 88.025 ;
        RECT 84.980 87.200 85.155 87.370 ;
        RECT 81.760 87.005 83.720 87.200 ;
        RECT 79.985 85.940 80.155 86.875 ;
        RECT 80.325 86.345 80.690 86.705 ;
        RECT 80.860 86.685 81.030 86.875 ;
        RECT 80.860 86.515 81.980 86.685 ;
        RECT 80.325 86.175 81.610 86.345 ;
        RECT 80.625 85.765 81.220 86.005 ;
        RECT 81.390 85.820 81.610 86.175 ;
        RECT 81.810 86.010 81.980 86.515 ;
        RECT 79.880 85.595 80.435 85.730 ;
        RECT 81.810 85.650 81.980 85.815 ;
        RECT 81.540 85.595 81.980 85.650 ;
        RECT 79.880 85.480 81.980 85.595 ;
        RECT 82.260 85.550 83.720 87.005 ;
        RECT 83.890 86.995 85.155 87.200 ;
        RECT 85.325 87.165 86.290 87.425 ;
        RECT 83.890 86.735 85.880 86.995 ;
        RECT 83.890 86.135 85.155 86.735 ;
        RECT 86.050 86.565 86.290 87.165 ;
        RECT 85.325 86.305 86.290 86.565 ;
        RECT 83.890 85.890 85.880 86.135 ;
        RECT 80.305 85.425 81.670 85.480 ;
        RECT 82.260 85.310 83.200 85.550 ;
        RECT 83.890 85.380 85.155 85.890 ;
        RECT 86.050 85.720 86.290 86.305 ;
        RECT 85.325 85.460 86.290 85.720 ;
        RECT 78.450 85.045 80.170 85.310 ;
        RECT 76.275 83.235 77.760 84.630 ;
        RECT 78.450 84.460 79.710 85.045 ;
        RECT 80.680 84.975 81.630 85.255 ;
        RECT 81.800 85.060 83.200 85.310 ;
        RECT 79.880 84.620 82.000 84.805 ;
        RECT 74.100 83.060 74.270 83.235 ;
        RECT 76.820 83.060 77.760 83.235 ;
        RECT 71.720 82.845 71.970 82.920 ;
        RECT 71.800 82.760 71.970 82.845 ;
        RECT 66.440 82.345 67.330 82.475 ;
        RECT 60.865 81.605 61.240 81.630 ;
        RECT 62.370 81.605 62.600 81.880 ;
        RECT 63.220 81.710 63.390 82.030 ;
        RECT 65.425 82.020 66.110 82.190 ;
        RECT 67.520 82.230 68.490 82.480 ;
        RECT 60.865 81.390 62.600 81.605 ;
        RECT 61.390 81.370 62.600 81.390 ;
        RECT 62.770 81.380 63.390 81.710 ;
        RECT 65.940 81.735 66.110 82.020 ;
        RECT 66.440 81.905 67.350 82.165 ;
        RECT 67.520 81.735 67.690 82.230 ;
        RECT 68.660 81.960 68.830 82.490 ;
        RECT 70.865 82.480 71.550 82.650 ;
        RECT 72.165 82.570 72.790 82.740 ;
        RECT 72.165 82.560 72.335 82.570 ;
        RECT 71.380 81.970 71.550 82.480 ;
        RECT 71.880 82.350 72.335 82.560 ;
        RECT 72.540 82.180 72.710 82.340 ;
        RECT 72.160 82.085 72.725 82.180 ;
        RECT 68.660 81.830 69.745 81.960 ;
        RECT 63.560 81.420 64.230 81.590 ;
        RECT 60.855 80.940 61.195 81.110 ;
        RECT 61.390 81.050 61.720 81.370 ;
        RECT 63.220 81.250 63.390 81.380 ;
        RECT 61.000 80.880 61.195 80.940 ;
        RECT 61.890 80.895 63.005 81.180 ;
        RECT 63.220 80.920 63.890 81.250 ;
        RECT 64.060 81.155 64.230 81.420 ;
        RECT 64.400 81.325 65.050 81.675 ;
        RECT 65.220 81.420 65.680 81.590 ;
        RECT 65.940 81.500 66.915 81.735 ;
        RECT 67.100 81.510 67.690 81.735 ;
        RECT 67.860 81.790 69.745 81.830 ;
        RECT 70.865 81.800 71.550 81.970 ;
        RECT 71.865 82.010 72.725 82.085 ;
        RECT 71.865 81.915 72.330 82.010 ;
        RECT 71.890 81.910 72.060 81.915 ;
        RECT 65.220 81.155 65.390 81.420 ;
        RECT 65.940 81.250 66.110 81.500 ;
        RECT 67.100 81.340 67.340 81.510 ;
        RECT 67.860 81.500 68.830 81.790 ;
        RECT 69.890 81.630 70.725 81.680 ;
        RECT 71.380 81.670 71.550 81.800 ;
        RECT 69.890 81.620 71.160 81.630 ;
        RECT 64.060 80.925 65.390 81.155 ;
        RECT 65.560 80.920 66.110 81.250 ;
        RECT 66.320 81.170 66.830 81.330 ;
        RECT 67.520 81.170 68.490 81.330 ;
        RECT 66.320 81.000 68.490 81.170 ;
        RECT 66.365 80.995 68.490 81.000 ;
        RECT 68.660 81.120 68.830 81.500 ;
        RECT 69.045 81.510 71.160 81.620 ;
        RECT 69.045 81.465 70.020 81.510 ;
        RECT 69.045 81.290 69.970 81.465 ;
        RECT 70.600 81.455 71.160 81.510 ;
        RECT 68.150 80.990 68.320 80.995 ;
        RECT 61.890 80.880 62.060 80.895 ;
        RECT 61.000 80.710 62.060 80.880 ;
        RECT 60.500 79.950 61.165 80.350 ;
        RECT 61.530 80.320 62.060 80.710 ;
        RECT 60.500 79.360 60.670 79.950 ;
        RECT 61.530 79.890 61.910 80.320 ;
        RECT 62.230 80.025 62.540 80.720 ;
        RECT 63.220 80.715 63.390 80.920 ;
        RECT 65.940 80.810 66.110 80.920 ;
        RECT 68.660 80.950 69.840 81.120 ;
        RECT 68.660 80.820 68.830 80.950 ;
        RECT 62.750 80.325 63.390 80.715 ;
        RECT 63.560 80.565 65.680 80.750 ;
        RECT 65.940 80.480 66.835 80.810 ;
        RECT 67.860 80.490 68.830 80.820 ;
        RECT 70.140 80.790 70.470 81.340 ;
        RECT 70.640 81.300 71.160 81.455 ;
        RECT 71.380 81.570 71.930 81.670 ;
        RECT 72.460 81.655 72.790 81.780 ;
        RECT 71.380 81.400 72.010 81.570 ;
        RECT 72.225 81.450 72.790 81.655 ;
        RECT 71.380 81.340 71.930 81.400 ;
        RECT 71.380 81.130 71.550 81.340 ;
        RECT 71.890 81.150 72.060 81.160 ;
        RECT 70.770 80.960 71.550 81.130 ;
        RECT 71.720 80.980 72.350 81.150 ;
        RECT 70.140 80.780 71.165 80.790 ;
        RECT 62.750 80.060 63.850 80.325 ;
        RECT 64.360 80.115 65.310 80.395 ;
        RECT 65.940 80.310 66.110 80.480 ;
        RECT 65.480 80.300 66.110 80.310 ;
        RECT 68.660 80.300 68.830 80.490 ;
        RECT 69.000 80.590 71.165 80.780 ;
        RECT 69.000 80.440 69.935 80.590 ;
        RECT 70.640 80.460 71.165 80.590 ;
        RECT 71.380 80.730 71.550 80.960 ;
        RECT 72.180 80.730 72.350 80.980 ;
        RECT 72.540 81.110 72.710 81.270 ;
        RECT 72.960 81.110 73.130 82.920 ;
        RECT 73.300 82.970 73.470 83.030 ;
        RECT 73.300 82.720 73.890 82.970 ;
        RECT 73.300 81.990 73.470 82.720 ;
        RECT 74.100 82.530 75.360 83.060 ;
        RECT 73.640 82.200 75.360 82.530 ;
        RECT 75.530 82.770 77.760 83.060 ;
        RECT 77.930 84.450 79.710 84.460 ;
        RECT 82.260 84.450 83.200 85.060 ;
        RECT 77.930 84.120 80.210 84.450 ;
        RECT 80.380 84.215 81.710 84.445 ;
        RECT 77.930 83.520 79.710 84.120 ;
        RECT 80.380 83.950 80.550 84.215 ;
        RECT 79.880 83.780 80.550 83.950 ;
        RECT 80.720 83.695 81.370 84.045 ;
        RECT 81.540 83.950 81.710 84.215 ;
        RECT 81.880 84.120 83.200 84.450 ;
        RECT 81.540 83.780 82.000 83.950 ;
        RECT 82.260 83.690 83.200 84.120 ;
        RECT 83.370 85.275 85.155 85.380 ;
        RECT 83.370 85.030 85.880 85.275 ;
        RECT 83.370 84.415 85.155 85.030 ;
        RECT 86.050 84.860 86.290 85.460 ;
        RECT 85.325 84.600 86.290 84.860 ;
        RECT 83.370 84.170 85.880 84.415 ;
        RECT 83.370 83.690 85.155 84.170 ;
        RECT 86.050 84.000 86.290 84.600 ;
        RECT 85.325 83.740 86.290 84.000 ;
        RECT 82.260 83.520 82.430 83.690 ;
        RECT 84.980 83.555 85.155 83.690 ;
        RECT 86.065 83.565 86.290 83.740 ;
        RECT 86.460 83.735 86.710 89.745 ;
        RECT 87.700 89.590 87.870 90.100 ;
        RECT 88.440 89.930 88.610 90.630 ;
        RECT 88.780 90.105 89.400 90.815 ;
        RECT 88.090 89.760 88.610 89.930 ;
        RECT 87.700 89.575 88.270 89.590 ;
        RECT 87.140 89.315 88.270 89.575 ;
        RECT 87.700 89.210 88.270 89.315 ;
        RECT 88.440 89.360 88.610 89.760 ;
        RECT 88.780 89.530 89.110 89.935 ;
        RECT 89.570 89.915 89.740 91.015 ;
        RECT 89.280 89.745 89.740 89.915 ;
        RECT 89.280 89.360 89.450 89.745 ;
        RECT 89.910 89.680 90.200 91.340 ;
        RECT 90.420 90.910 91.430 91.340 ;
        RECT 91.600 90.950 92.920 91.340 ;
        RECT 90.420 90.320 90.590 90.910 ;
        RECT 91.600 90.740 91.810 90.950 ;
        RECT 91.100 90.490 91.810 90.740 ;
        RECT 90.420 90.070 91.090 90.320 ;
        RECT 90.420 89.510 90.590 90.070 ;
        RECT 86.880 88.885 87.505 89.145 ;
        RECT 86.880 88.285 87.050 88.885 ;
        RECT 87.700 88.715 87.870 89.210 ;
        RECT 88.440 89.190 89.450 89.360 ;
        RECT 89.620 89.230 90.590 89.510 ;
        RECT 88.780 89.085 89.110 89.190 ;
        RECT 88.200 88.915 88.545 89.020 ;
        RECT 89.280 88.915 90.250 89.020 ;
        RECT 88.200 88.745 90.250 88.915 ;
        RECT 87.220 88.575 87.870 88.715 ;
        RECT 90.420 88.575 90.590 89.230 ;
        RECT 90.760 89.550 91.090 89.800 ;
        RECT 90.760 89.000 90.930 89.550 ;
        RECT 91.260 89.380 91.430 90.490 ;
        RECT 91.980 90.250 92.150 90.740 ;
        RECT 91.100 89.170 91.430 89.380 ;
        RECT 91.600 90.080 92.150 90.250 ;
        RECT 92.320 90.450 92.580 90.780 ;
        RECT 90.760 88.675 91.100 89.000 ;
        RECT 91.600 88.925 91.770 90.080 ;
        RECT 92.320 89.420 92.500 90.450 ;
        RECT 92.750 90.030 92.920 90.950 ;
        RECT 93.140 91.175 93.310 91.510 ;
        RECT 93.505 91.345 94.130 91.605 ;
        RECT 93.140 90.915 93.790 91.175 ;
        RECT 93.140 90.315 93.310 90.915 ;
        RECT 93.960 90.745 94.130 91.345 ;
        RECT 93.505 90.485 94.130 90.745 ;
        RECT 93.140 90.055 93.870 90.315 ;
        RECT 93.140 89.760 93.310 90.055 ;
        RECT 94.300 89.885 94.550 95.895 ;
        RECT 94.720 95.890 94.945 96.065 ;
        RECT 94.720 95.630 95.685 95.890 ;
        RECT 94.720 95.030 94.960 95.630 ;
        RECT 95.855 95.460 96.030 96.075 ;
        RECT 95.130 95.215 96.030 95.460 ;
        RECT 94.720 94.770 95.685 95.030 ;
        RECT 94.720 94.170 94.960 94.770 ;
        RECT 95.855 94.600 96.030 95.215 ;
        RECT 96.200 95.770 96.880 96.540 ;
        RECT 97.050 96.010 97.220 98.405 ;
        RECT 97.390 97.395 97.590 98.745 ;
        RECT 98.110 98.690 98.750 98.755 ;
        RECT 98.110 98.585 99.570 98.690 ;
        RECT 98.580 98.415 99.570 98.585 ;
        RECT 99.740 98.415 99.940 99.135 ;
        RECT 100.120 98.690 100.330 99.360 ;
        RECT 101.300 99.190 102.560 99.620 ;
        RECT 100.500 98.860 102.560 99.190 ;
        RECT 102.730 99.485 104.660 99.620 ;
        RECT 102.730 98.870 104.190 99.485 ;
        RECT 104.830 99.315 105.010 99.825 ;
        RECT 104.360 98.950 105.010 99.315 ;
        RECT 105.180 99.825 105.720 99.995 ;
        RECT 105.890 101.935 106.070 102.525 ;
        RECT 106.740 102.355 106.910 103.010 ;
        RECT 106.240 102.105 106.910 102.355 ;
        RECT 107.080 103.240 107.410 103.315 ;
        RECT 107.080 103.070 107.420 103.240 ;
        RECT 107.080 103.065 107.410 103.070 ;
        RECT 107.080 102.475 107.250 103.065 ;
        RECT 107.590 102.895 107.760 104.015 ;
        RECT 108.640 103.775 108.820 104.015 ;
        RECT 108.990 103.945 110.175 104.115 ;
        RECT 108.270 103.600 108.470 103.760 ;
        RECT 107.420 102.645 107.760 102.895 ;
        RECT 107.080 102.225 107.410 102.475 ;
        RECT 107.590 102.255 107.760 102.645 ;
        RECT 107.930 103.430 108.470 103.600 ;
        RECT 108.640 103.445 109.290 103.775 ;
        RECT 107.930 102.595 108.100 103.430 ;
        RECT 108.270 102.765 108.470 103.260 ;
        RECT 108.640 102.935 108.820 103.445 ;
        RECT 109.460 103.275 110.175 103.945 ;
        RECT 108.990 103.105 110.175 103.275 ;
        RECT 108.640 102.605 109.290 102.935 ;
        RECT 109.460 102.635 110.175 103.105 ;
        RECT 107.930 102.425 108.470 102.595 ;
        RECT 109.460 102.435 111.005 102.635 ;
        RECT 105.890 101.685 106.570 101.935 ;
        RECT 105.890 101.095 106.070 101.685 ;
        RECT 106.740 101.535 106.910 102.105 ;
        RECT 107.590 102.085 108.100 102.255 ;
        RECT 107.080 101.915 107.420 102.020 ;
        RECT 107.080 101.705 107.760 101.915 ;
        RECT 106.740 101.515 107.410 101.535 ;
        RECT 106.240 101.285 107.410 101.515 ;
        RECT 106.240 101.265 106.910 101.285 ;
        RECT 105.890 100.845 106.570 101.095 ;
        RECT 105.180 98.970 105.390 99.825 ;
        RECT 105.890 99.615 106.060 100.845 ;
        RECT 106.740 100.695 106.910 101.265 ;
        RECT 107.590 101.115 107.760 101.705 ;
        RECT 107.080 100.865 107.760 101.115 ;
        RECT 106.230 100.285 106.570 100.535 ;
        RECT 106.740 100.390 107.410 100.695 ;
        RECT 106.740 100.115 106.910 100.390 ;
        RECT 107.590 100.220 107.760 100.865 ;
        RECT 106.240 99.865 106.910 100.115 ;
        RECT 105.560 99.445 106.060 99.615 ;
        RECT 101.300 98.700 102.560 98.860 ;
        RECT 103.250 98.780 104.190 98.870 ;
        RECT 100.120 98.415 101.130 98.690 ;
        RECT 97.760 97.985 98.410 98.315 ;
        RECT 98.580 98.240 98.750 98.415 ;
        RECT 101.300 98.240 103.080 98.700 ;
        RECT 97.760 97.475 97.940 97.985 ;
        RECT 98.580 97.815 100.040 98.240 ;
        RECT 98.110 97.645 100.040 97.815 ;
        RECT 98.580 97.490 100.040 97.645 ;
        RECT 100.210 97.950 103.080 98.240 ;
        RECT 103.250 98.610 104.660 98.780 ;
        RECT 103.250 97.950 104.190 98.610 ;
        RECT 97.760 97.225 98.410 97.475 ;
        RECT 97.390 96.535 97.590 97.205 ;
        RECT 97.760 96.670 98.020 97.000 ;
        RECT 97.050 95.840 97.590 96.010 ;
        RECT 96.200 95.180 96.370 95.770 ;
        RECT 96.540 95.350 97.250 95.600 ;
        RECT 97.420 95.350 97.590 95.840 ;
        RECT 97.760 95.640 97.940 96.670 ;
        RECT 98.190 96.245 98.410 97.225 ;
        RECT 98.580 96.570 99.520 97.490 ;
        RECT 100.210 97.320 101.470 97.950 ;
        RECT 101.640 97.550 103.460 97.780 ;
        RECT 101.640 97.465 102.320 97.550 ;
        RECT 99.690 97.295 101.470 97.320 ;
        RECT 99.690 97.045 101.970 97.295 ;
        RECT 99.690 96.570 101.470 97.045 ;
        RECT 102.140 96.875 102.320 97.465 ;
        RECT 102.820 97.075 103.030 97.380 ;
        RECT 101.640 96.625 102.320 96.875 ;
        RECT 98.580 96.400 98.750 96.570 ;
        RECT 101.300 96.455 101.470 96.570 ;
        RECT 101.300 96.400 101.970 96.455 ;
        RECT 98.580 96.125 99.410 96.400 ;
        RECT 98.580 95.980 98.750 96.125 ;
        RECT 98.110 95.810 98.750 95.980 ;
        RECT 99.590 95.970 100.110 96.400 ;
        RECT 100.290 96.205 101.970 96.400 ;
        RECT 100.290 96.140 101.470 96.205 ;
        RECT 99.590 95.955 101.130 95.970 ;
        RECT 96.200 94.930 96.870 95.180 ;
        RECT 97.040 95.140 97.250 95.350 ;
        RECT 97.760 95.310 98.020 95.640 ;
        RECT 98.580 95.530 98.750 95.810 ;
        RECT 98.920 95.800 101.130 95.955 ;
        RECT 98.920 95.785 100.110 95.800 ;
        RECT 98.920 95.705 99.380 95.785 ;
        RECT 100.460 95.695 101.130 95.800 ;
        RECT 97.760 95.140 97.940 95.310 ;
        RECT 98.580 95.200 99.245 95.530 ;
        RECT 99.660 95.385 100.260 95.615 ;
        RECT 101.300 95.495 101.470 96.140 ;
        RECT 102.140 96.035 102.320 96.625 ;
        RECT 101.640 95.785 102.320 96.035 ;
        RECT 98.580 95.140 98.750 95.200 ;
        RECT 97.040 94.730 97.940 95.140 ;
        RECT 98.110 94.970 98.750 95.140 ;
        RECT 99.415 95.020 99.910 95.200 ;
        RECT 95.130 94.355 96.030 94.600 ;
        RECT 94.720 93.910 95.685 94.170 ;
        RECT 95.855 94.080 96.030 94.355 ;
        RECT 96.200 94.390 98.410 94.560 ;
        RECT 96.200 94.250 97.170 94.390 ;
        RECT 98.080 94.260 98.410 94.390 ;
        RECT 94.720 93.325 94.960 93.910 ;
        RECT 95.855 93.770 96.830 94.080 ;
        RECT 95.855 93.740 96.030 93.770 ;
        RECT 95.130 93.495 96.030 93.740 ;
        RECT 97.000 93.700 97.170 94.250 ;
        RECT 97.340 93.870 97.910 94.220 ;
        RECT 98.580 94.090 98.750 94.970 ;
        RECT 98.970 94.790 99.910 95.020 ;
        RECT 100.090 95.055 100.260 95.385 ;
        RECT 100.455 95.280 101.470 95.495 ;
        RECT 100.090 94.805 100.555 95.055 ;
        RECT 100.090 94.620 100.260 94.805 ;
        RECT 100.790 94.620 101.130 95.095 ;
        RECT 101.300 95.055 101.470 95.280 ;
        RECT 101.640 95.225 101.980 95.475 ;
        RECT 101.300 94.805 101.970 95.055 ;
        RECT 98.100 93.815 98.750 94.090 ;
        RECT 98.970 94.365 100.260 94.620 ;
        RECT 98.970 93.830 99.235 94.365 ;
        RECT 94.720 93.065 95.685 93.325 ;
        RECT 95.855 93.170 96.030 93.495 ;
        RECT 96.200 93.340 96.830 93.600 ;
        RECT 97.000 93.530 97.590 93.700 ;
        RECT 98.580 93.640 98.750 93.815 ;
        RECT 99.430 93.810 99.910 94.195 ;
        RECT 100.090 94.080 100.260 94.365 ;
        RECT 100.430 94.440 100.620 94.580 ;
        RECT 101.300 94.440 101.470 94.805 ;
        RECT 100.430 94.250 101.470 94.440 ;
        RECT 100.090 93.825 100.625 94.080 ;
        RECT 100.795 93.810 101.470 94.250 ;
        RECT 101.300 93.640 101.470 93.810 ;
        RECT 94.720 92.465 94.960 93.065 ;
        RECT 95.855 92.915 96.490 93.170 ;
        RECT 95.855 92.895 96.030 92.915 ;
        RECT 95.130 92.635 96.030 92.895 ;
        RECT 96.660 92.740 96.830 93.340 ;
        RECT 94.720 92.205 95.685 92.465 ;
        RECT 95.855 92.310 96.030 92.635 ;
        RECT 96.200 92.480 97.250 92.740 ;
        RECT 97.420 92.560 97.590 93.530 ;
        RECT 97.760 93.340 98.320 93.635 ;
        RECT 97.760 92.740 97.930 93.340 ;
        RECT 98.580 93.170 99.295 93.640 ;
        RECT 98.100 92.915 99.295 93.170 ;
        RECT 97.080 92.390 97.250 92.480 ;
        RECT 97.760 92.480 98.320 92.740 ;
        RECT 97.760 92.390 97.930 92.480 ;
        RECT 94.720 91.605 94.960 92.205 ;
        RECT 95.855 92.035 96.900 92.310 ;
        RECT 95.130 92.025 96.900 92.035 ;
        RECT 95.130 91.800 96.030 92.025 ;
        RECT 97.080 91.985 97.930 92.390 ;
        RECT 98.580 92.310 99.295 92.915 ;
        RECT 98.100 92.055 99.295 92.310 ;
        RECT 100.865 93.240 101.470 93.640 ;
        RECT 101.640 94.310 101.980 94.635 ;
        RECT 102.150 94.555 102.320 95.785 ;
        RECT 102.490 96.905 103.030 97.075 ;
        RECT 103.210 97.005 103.460 97.550 ;
        RECT 102.490 94.935 102.660 96.905 ;
        RECT 103.630 96.835 103.850 97.760 ;
        RECT 102.830 95.160 103.030 96.610 ;
        RECT 103.200 96.585 103.850 96.835 ;
        RECT 103.200 96.075 103.380 96.585 ;
        RECT 104.020 96.415 104.190 97.950 ;
        RECT 104.410 97.420 104.580 98.340 ;
        RECT 104.830 97.920 105.010 98.950 ;
        RECT 105.560 98.290 105.730 99.445 ;
        RECT 106.230 99.370 106.570 99.695 ;
        RECT 104.750 97.590 105.010 97.920 ;
        RECT 105.180 98.120 105.730 98.290 ;
        RECT 105.900 98.990 106.230 99.200 ;
        RECT 105.180 97.630 105.350 98.120 ;
        RECT 105.900 97.880 106.070 98.990 ;
        RECT 106.400 98.820 106.570 99.370 ;
        RECT 106.240 98.570 106.570 98.820 ;
        RECT 106.740 98.300 106.910 99.865 ;
        RECT 107.080 99.450 107.760 100.220 ;
        RECT 107.930 99.690 108.100 102.085 ;
        RECT 108.270 101.075 108.470 102.425 ;
        RECT 108.990 102.295 111.005 102.435 ;
        RECT 108.990 102.265 110.175 102.295 ;
        RECT 108.640 101.665 109.290 101.995 ;
        RECT 108.640 101.155 108.820 101.665 ;
        RECT 109.460 101.495 110.175 102.265 ;
        RECT 108.990 101.325 110.175 101.495 ;
        RECT 108.640 100.905 109.290 101.155 ;
        RECT 108.270 100.215 108.470 100.885 ;
        RECT 108.640 100.350 108.900 100.680 ;
        RECT 107.930 99.520 108.470 99.690 ;
        RECT 107.080 98.860 107.250 99.450 ;
        RECT 107.420 99.030 108.130 99.280 ;
        RECT 108.300 99.030 108.470 99.520 ;
        RECT 108.640 99.320 108.820 100.350 ;
        RECT 109.070 99.925 109.290 100.905 ;
        RECT 109.460 99.660 110.175 101.325 ;
        RECT 111.745 100.815 112.350 104.220 ;
        RECT 110.495 100.465 112.350 100.815 ;
        RECT 108.990 99.490 110.175 99.660 ;
        RECT 107.080 98.610 107.750 98.860 ;
        RECT 107.920 98.820 108.130 99.030 ;
        RECT 108.640 98.990 108.900 99.320 ;
        RECT 108.640 98.820 108.820 98.990 ;
        RECT 109.460 98.875 110.175 99.490 ;
        RECT 111.745 98.875 112.350 100.465 ;
        RECT 109.460 98.820 109.630 98.875 ;
        RECT 107.920 98.410 108.820 98.820 ;
        RECT 108.990 98.700 109.630 98.820 ;
        RECT 112.180 98.700 112.350 98.875 ;
        RECT 108.990 98.650 110.175 98.700 ;
        RECT 106.240 98.050 106.910 98.300 ;
        RECT 105.520 97.630 106.230 97.880 ;
        RECT 106.740 97.755 106.910 98.050 ;
        RECT 107.080 98.010 108.900 98.240 ;
        RECT 107.080 97.925 107.760 98.010 ;
        RECT 105.520 97.420 105.730 97.630 ;
        RECT 106.740 97.505 107.410 97.755 ;
        RECT 106.740 97.460 106.910 97.505 ;
        RECT 104.410 97.030 105.730 97.420 ;
        RECT 105.900 97.030 106.910 97.460 ;
        RECT 107.580 97.335 107.760 97.925 ;
        RECT 108.260 97.535 108.470 97.840 ;
        RECT 107.080 97.085 107.760 97.335 ;
        RECT 103.550 96.245 104.190 96.415 ;
        RECT 104.020 96.230 104.190 96.245 ;
        RECT 106.740 96.915 106.910 97.030 ;
        RECT 106.740 96.665 107.410 96.915 ;
        RECT 103.200 95.745 103.850 96.075 ;
        RECT 104.020 96.060 104.705 96.230 ;
        RECT 106.740 96.220 106.910 96.665 ;
        RECT 107.580 96.495 107.760 97.085 ;
        RECT 107.080 96.245 107.760 96.495 ;
        RECT 104.020 95.435 104.190 96.060 ;
        RECT 105.825 96.050 106.910 96.220 ;
        RECT 104.845 95.890 105.680 95.940 ;
        RECT 104.410 95.880 105.680 95.890 ;
        RECT 104.410 95.770 106.525 95.880 ;
        RECT 104.410 95.715 104.970 95.770 ;
        RECT 105.550 95.725 106.525 95.770 ;
        RECT 104.410 95.560 104.930 95.715 ;
        RECT 103.200 95.390 104.190 95.435 ;
        RECT 103.200 95.265 104.800 95.390 ;
        RECT 104.020 95.220 104.800 95.265 ;
        RECT 102.490 94.765 103.030 94.935 ;
        RECT 102.150 94.385 102.650 94.555 ;
        RECT 101.640 93.760 101.810 94.310 ;
        RECT 101.980 93.930 102.310 94.140 ;
        RECT 101.640 93.510 101.970 93.760 ;
        RECT 100.865 92.990 101.970 93.240 ;
        RECT 100.865 92.400 101.470 92.990 ;
        RECT 102.140 92.820 102.310 93.930 ;
        RECT 102.480 93.230 102.650 94.385 ;
        RECT 102.820 93.910 103.030 94.765 ;
        RECT 103.200 94.765 103.850 95.095 ;
        RECT 103.200 94.255 103.380 94.765 ;
        RECT 104.020 94.595 104.190 95.220 ;
        RECT 105.100 95.050 105.430 95.600 ;
        RECT 105.600 95.550 106.525 95.725 ;
        RECT 106.740 95.515 106.910 96.050 ;
        RECT 107.080 95.685 107.420 95.935 ;
        RECT 106.740 95.380 107.410 95.515 ;
        RECT 105.730 95.265 107.410 95.380 ;
        RECT 105.730 95.210 106.910 95.265 ;
        RECT 104.405 95.040 105.430 95.050 ;
        RECT 104.405 94.850 106.570 95.040 ;
        RECT 104.405 94.720 104.930 94.850 ;
        RECT 105.635 94.700 106.570 94.850 ;
        RECT 103.550 94.460 104.190 94.595 ;
        RECT 103.550 94.425 104.720 94.460 ;
        RECT 103.200 93.890 103.850 94.255 ;
        RECT 104.020 94.250 104.720 94.425 ;
        RECT 102.480 93.060 103.030 93.230 ;
        RECT 101.980 92.570 102.690 92.820 ;
        RECT 102.860 92.570 103.030 93.060 ;
        RECT 103.200 92.860 103.380 93.890 ;
        RECT 104.020 93.720 104.190 94.250 ;
        RECT 105.100 93.975 105.430 94.680 ;
        RECT 105.635 94.145 106.010 94.700 ;
        RECT 106.740 94.470 106.910 95.210 ;
        RECT 106.240 94.155 106.910 94.470 ;
        RECT 103.550 93.550 104.190 93.720 ;
        RECT 98.100 92.030 100.125 92.055 ;
        RECT 98.580 91.800 100.125 92.030 ;
        RECT 95.130 91.775 97.195 91.800 ;
        RECT 94.720 91.345 95.685 91.605 ;
        RECT 95.855 91.510 97.195 91.775 ;
        RECT 97.855 91.715 100.125 91.800 ;
        RECT 100.865 91.970 102.310 92.400 ;
        RECT 102.480 92.360 102.690 92.570 ;
        RECT 103.200 92.530 103.460 92.860 ;
        RECT 103.630 92.360 103.800 93.280 ;
        RECT 102.480 91.970 103.800 92.360 ;
        RECT 104.020 92.435 104.190 93.550 ;
        RECT 104.470 93.805 106.440 93.975 ;
        RECT 104.470 93.190 104.640 93.805 ;
        RECT 104.810 93.315 106.100 93.635 ;
        RECT 104.810 93.170 105.140 93.315 ;
        RECT 104.470 92.785 104.640 93.020 ;
        RECT 105.350 92.955 106.070 93.145 ;
        RECT 106.270 93.090 106.440 93.805 ;
        RECT 106.740 93.700 106.910 94.155 ;
        RECT 107.080 94.770 107.420 95.095 ;
        RECT 107.590 95.015 107.760 96.245 ;
        RECT 107.930 97.365 108.470 97.535 ;
        RECT 108.650 97.465 108.900 98.010 ;
        RECT 107.930 95.395 108.100 97.365 ;
        RECT 109.070 97.295 109.290 98.220 ;
        RECT 108.270 95.620 108.470 97.070 ;
        RECT 108.640 97.045 109.290 97.295 ;
        RECT 109.460 97.115 110.175 98.650 ;
        RECT 108.640 96.535 108.820 97.045 ;
        RECT 109.460 96.875 111.005 97.115 ;
        RECT 108.990 96.775 111.005 96.875 ;
        RECT 108.990 96.705 110.175 96.775 ;
        RECT 108.640 96.205 109.290 96.535 ;
        RECT 109.460 95.895 110.175 96.705 ;
        RECT 108.640 95.725 110.175 95.895 ;
        RECT 107.930 95.225 108.470 95.395 ;
        RECT 107.590 94.845 108.090 95.015 ;
        RECT 107.080 94.220 107.250 94.770 ;
        RECT 107.420 94.390 107.750 94.600 ;
        RECT 107.080 93.970 107.410 94.220 ;
        RECT 106.740 93.450 107.410 93.700 ;
        RECT 106.240 92.785 106.570 92.865 ;
        RECT 104.470 92.615 106.570 92.785 ;
        RECT 106.740 92.860 106.910 93.450 ;
        RECT 107.580 93.280 107.750 94.390 ;
        RECT 107.920 93.690 108.090 94.845 ;
        RECT 108.260 94.370 108.470 95.225 ;
        RECT 108.640 95.225 109.290 95.555 ;
        RECT 108.640 94.715 108.820 95.225 ;
        RECT 109.460 95.055 110.175 95.725 ;
        RECT 111.745 95.295 112.350 98.700 ;
        RECT 108.990 94.885 110.175 95.055 ;
        RECT 110.495 94.945 112.350 95.295 ;
        RECT 108.640 94.350 109.290 94.715 ;
        RECT 107.920 93.520 108.470 93.690 ;
        RECT 107.420 93.030 108.130 93.280 ;
        RECT 108.300 93.030 108.470 93.520 ;
        RECT 108.640 93.320 108.820 94.350 ;
        RECT 109.460 94.180 110.175 94.885 ;
        RECT 108.990 94.010 110.175 94.180 ;
        RECT 104.020 92.065 104.690 92.435 ;
        RECT 104.870 92.155 105.170 92.615 ;
        RECT 106.740 92.445 107.750 92.860 ;
        RECT 105.350 92.275 105.680 92.445 ;
        RECT 105.940 92.430 107.750 92.445 ;
        RECT 107.920 92.820 108.130 93.030 ;
        RECT 108.640 92.990 108.900 93.320 ;
        RECT 109.070 92.820 109.240 93.740 ;
        RECT 107.920 92.430 109.240 92.820 ;
        RECT 109.460 93.355 110.175 94.010 ;
        RECT 111.745 93.355 112.350 94.945 ;
        RECT 109.460 93.180 109.630 93.355 ;
        RECT 112.180 93.180 112.350 93.355 ;
        RECT 109.460 92.660 110.920 93.180 ;
        RECT 105.940 92.275 106.910 92.430 ;
        RECT 100.865 91.800 101.470 91.970 ;
        RECT 104.020 91.800 104.190 92.065 ;
        RECT 104.870 91.955 105.200 92.155 ;
        RECT 105.420 92.105 105.680 92.275 ;
        RECT 97.855 91.510 99.295 91.715 ;
        RECT 94.720 90.745 94.960 91.345 ;
        RECT 95.855 91.175 96.030 91.510 ;
        RECT 95.130 90.915 96.030 91.175 ;
        RECT 94.720 90.485 95.685 90.745 ;
        RECT 95.855 90.315 96.030 90.915 ;
        RECT 95.060 90.055 96.030 90.315 ;
        RECT 96.200 91.000 96.830 91.300 ;
        RECT 98.580 91.290 99.295 91.510 ;
        RECT 97.050 91.260 97.220 91.280 ;
        RECT 97.000 91.045 97.930 91.260 ;
        RECT 96.200 90.330 96.370 91.000 ;
        RECT 97.000 90.830 97.220 91.045 ;
        RECT 96.540 90.500 97.220 90.830 ;
        RECT 96.200 90.160 97.210 90.330 ;
        RECT 95.860 89.990 96.030 90.055 ;
        RECT 92.670 89.590 93.310 89.760 ;
        RECT 93.490 89.635 95.685 89.885 ;
        RECT 95.860 89.660 96.830 89.990 ;
        RECT 93.140 89.455 93.310 89.590 ;
        RECT 91.270 88.755 91.770 88.925 ;
        RECT 87.220 88.455 88.785 88.575 ;
        RECT 87.700 88.405 88.785 88.455 ;
        RECT 89.240 88.505 90.590 88.575 ;
        RECT 89.240 88.405 91.090 88.505 ;
        RECT 86.880 88.025 87.505 88.285 ;
        RECT 87.700 88.120 87.870 88.405 ;
        RECT 90.420 88.255 91.090 88.405 ;
        RECT 90.420 88.120 90.590 88.255 ;
        RECT 86.880 87.425 87.050 88.025 ;
        RECT 87.700 87.855 88.415 88.120 ;
        RECT 87.220 87.595 88.415 87.855 ;
        RECT 86.880 87.165 87.505 87.425 ;
        RECT 86.880 86.580 87.050 87.165 ;
        RECT 87.700 86.995 88.415 87.595 ;
        RECT 87.220 86.750 88.415 86.995 ;
        RECT 86.880 86.305 87.505 86.580 ;
        RECT 87.700 86.535 88.415 86.750 ;
        RECT 89.985 87.105 90.590 88.120 ;
        RECT 90.760 87.835 91.100 88.085 ;
        RECT 91.270 87.525 91.440 88.755 ;
        RECT 91.940 88.545 92.150 89.400 ;
        RECT 90.760 87.275 91.440 87.525 ;
        RECT 89.985 86.855 91.090 87.105 ;
        RECT 86.880 85.720 87.050 86.305 ;
        RECT 87.700 86.195 89.245 86.535 ;
        RECT 89.985 86.265 90.590 86.855 ;
        RECT 91.260 86.685 91.440 87.275 ;
        RECT 90.760 86.435 91.440 86.685 ;
        RECT 87.700 86.135 88.415 86.195 ;
        RECT 87.220 85.890 88.415 86.135 ;
        RECT 86.880 85.460 87.505 85.720 ;
        RECT 86.880 84.860 87.050 85.460 ;
        RECT 87.700 85.280 88.415 85.890 ;
        RECT 87.220 85.030 88.415 85.280 ;
        RECT 86.880 84.600 87.505 84.860 ;
        RECT 86.880 84.000 87.050 84.600 ;
        RECT 87.700 84.420 88.415 85.030 ;
        RECT 89.985 86.015 91.090 86.265 ;
        RECT 89.985 85.360 90.590 86.015 ;
        RECT 91.260 85.845 91.440 86.435 ;
        RECT 91.610 88.375 92.150 88.545 ;
        RECT 92.320 89.055 92.970 89.420 ;
        RECT 93.140 89.195 93.835 89.455 ;
        RECT 92.320 88.545 92.500 89.055 ;
        RECT 93.140 88.885 93.310 89.195 ;
        RECT 94.300 89.025 94.550 89.635 ;
        RECT 95.860 89.455 96.030 89.660 ;
        RECT 97.000 89.490 97.210 90.160 ;
        RECT 97.390 90.105 97.590 90.875 ;
        RECT 97.760 90.830 97.930 91.045 ;
        RECT 98.110 91.000 99.295 91.290 ;
        RECT 97.760 90.500 98.410 90.830 ;
        RECT 97.760 89.990 97.940 90.500 ;
        RECT 98.580 90.330 99.295 91.000 ;
        RECT 98.110 90.160 99.295 90.330 ;
        RECT 100.865 91.510 102.635 91.800 ;
        RECT 103.295 91.510 104.190 91.800 ;
        RECT 105.420 91.935 106.465 92.105 ;
        RECT 105.420 91.745 105.590 91.935 ;
        RECT 100.865 91.340 101.470 91.510 ;
        RECT 100.865 90.910 102.310 91.340 ;
        RECT 102.480 90.950 103.800 91.340 ;
        RECT 100.865 90.320 101.470 90.910 ;
        RECT 102.480 90.740 102.690 90.950 ;
        RECT 101.980 90.490 102.690 90.740 ;
        RECT 100.865 90.235 101.970 90.320 ;
        RECT 95.050 89.195 96.030 89.455 ;
        RECT 96.200 89.215 97.210 89.490 ;
        RECT 97.390 89.215 97.590 89.935 ;
        RECT 97.760 89.660 98.410 89.990 ;
        RECT 98.580 89.490 99.295 90.160 ;
        RECT 99.615 90.070 101.970 90.235 ;
        RECT 99.615 89.885 101.470 90.070 ;
        RECT 97.760 89.215 99.295 89.490 ;
        RECT 92.670 88.715 93.310 88.885 ;
        RECT 93.490 89.020 94.550 89.025 ;
        RECT 95.860 89.040 96.030 89.195 ;
        RECT 98.580 89.040 99.295 89.215 ;
        RECT 93.490 88.775 95.690 89.020 ;
        RECT 93.140 88.595 93.310 88.715 ;
        RECT 91.610 86.405 91.780 88.375 ;
        RECT 92.320 88.215 92.970 88.545 ;
        RECT 93.140 88.290 93.820 88.595 ;
        RECT 93.990 88.290 94.550 88.605 ;
        RECT 95.860 88.595 97.120 89.040 ;
        RECT 95.050 88.300 97.120 88.595 ;
        RECT 91.950 86.700 92.150 88.150 ;
        RECT 93.140 88.045 93.310 88.290 ;
        RECT 92.320 87.950 93.310 88.045 ;
        RECT 92.320 87.875 93.825 87.950 ;
        RECT 95.860 87.940 97.120 88.300 ;
        RECT 93.140 87.780 93.825 87.875 ;
        RECT 92.320 87.235 92.970 87.565 ;
        RECT 92.320 86.725 92.500 87.235 ;
        RECT 93.140 87.110 93.310 87.780 ;
        RECT 94.945 87.770 97.120 87.940 ;
        RECT 97.290 88.295 99.295 89.040 ;
        RECT 100.865 88.505 101.470 89.885 ;
        RECT 101.640 89.550 101.970 89.800 ;
        RECT 101.640 89.000 101.810 89.550 ;
        RECT 102.140 89.380 102.310 90.490 ;
        RECT 102.860 90.250 103.030 90.740 ;
        RECT 101.980 89.170 102.310 89.380 ;
        RECT 102.480 90.080 103.030 90.250 ;
        RECT 103.200 90.450 103.460 90.780 ;
        RECT 101.640 88.675 101.980 89.000 ;
        RECT 102.480 88.925 102.650 90.080 ;
        RECT 103.200 89.420 103.380 90.450 ;
        RECT 103.630 90.030 103.800 90.950 ;
        RECT 104.020 90.370 104.190 91.510 ;
        RECT 104.470 91.575 105.590 91.745 ;
        RECT 104.470 91.070 104.640 91.575 ;
        RECT 105.760 91.405 106.125 91.765 ;
        RECT 104.840 91.235 106.125 91.405 ;
        RECT 104.840 90.880 105.060 91.235 ;
        RECT 104.470 90.710 104.640 90.875 ;
        RECT 105.230 90.825 105.825 91.065 ;
        RECT 106.295 91.000 106.465 91.935 ;
        RECT 106.740 91.800 106.910 92.275 ;
        RECT 109.460 91.970 110.380 92.660 ;
        RECT 111.090 92.490 112.350 93.180 ;
        RECT 110.550 91.970 112.350 92.490 ;
        RECT 109.460 91.800 109.630 91.970 ;
        RECT 112.180 91.800 112.350 91.970 ;
        RECT 106.740 91.510 108.075 91.800 ;
        RECT 108.735 91.510 110.355 91.800 ;
        RECT 111.015 91.510 112.350 91.800 ;
        RECT 104.470 90.655 104.910 90.710 ;
        RECT 106.015 90.655 106.570 90.790 ;
        RECT 104.470 90.540 106.570 90.655 ;
        RECT 104.780 90.485 106.145 90.540 ;
        RECT 106.740 90.420 106.910 91.510 ;
        RECT 109.460 91.340 109.630 91.510 ;
        RECT 112.180 91.340 112.350 91.510 ;
        RECT 109.460 90.420 110.175 91.340 ;
        RECT 106.740 90.370 108.050 90.420 ;
        RECT 104.020 90.120 104.650 90.370 ;
        RECT 104.020 89.760 104.190 90.120 ;
        RECT 104.820 90.035 105.770 90.315 ;
        RECT 106.280 90.130 108.050 90.370 ;
        RECT 108.660 90.130 110.175 90.420 ;
        RECT 106.280 90.105 106.910 90.130 ;
        RECT 103.550 89.590 104.190 89.760 ;
        RECT 104.450 89.680 106.570 89.865 ;
        RECT 104.020 89.510 104.190 89.590 ;
        RECT 106.740 89.510 106.910 90.105 ;
        RECT 107.080 89.710 109.290 89.960 ;
        RECT 107.080 89.510 107.630 89.710 ;
        RECT 102.150 88.755 102.650 88.925 ;
        RECT 100.865 88.295 101.970 88.505 ;
        RECT 97.290 88.120 98.750 88.295 ;
        RECT 101.300 88.255 101.970 88.295 ;
        RECT 101.300 88.120 101.470 88.255 ;
        RECT 97.290 87.830 99.295 88.120 ;
        RECT 95.860 87.660 97.120 87.770 ;
        RECT 93.965 87.610 94.800 87.660 ;
        RECT 93.530 87.600 94.800 87.610 ;
        RECT 93.530 87.490 95.645 87.600 ;
        RECT 93.530 87.435 94.090 87.490 ;
        RECT 94.670 87.445 95.645 87.490 ;
        RECT 93.530 87.280 94.050 87.435 ;
        RECT 93.140 87.065 93.920 87.110 ;
        RECT 92.670 86.940 93.920 87.065 ;
        RECT 92.670 86.895 93.310 86.940 ;
        RECT 92.320 86.475 92.970 86.725 ;
        RECT 91.610 86.235 92.150 86.405 ;
        RECT 91.940 85.930 92.150 86.235 ;
        RECT 90.760 85.760 91.440 85.845 ;
        RECT 92.330 85.760 92.580 86.305 ;
        RECT 90.760 85.530 92.580 85.760 ;
        RECT 92.750 85.550 92.970 86.475 ;
        RECT 93.140 86.180 93.310 86.895 ;
        RECT 94.220 86.770 94.550 87.320 ;
        RECT 94.720 87.270 95.645 87.445 ;
        RECT 95.860 87.100 97.640 87.660 ;
        RECT 94.850 86.930 97.640 87.100 ;
        RECT 93.525 86.760 94.550 86.770 ;
        RECT 93.525 86.570 95.690 86.760 ;
        RECT 93.525 86.440 94.050 86.570 ;
        RECT 94.755 86.420 95.690 86.570 ;
        RECT 95.860 86.450 97.640 86.930 ;
        RECT 97.810 86.535 99.295 87.830 ;
        RECT 100.865 87.105 101.470 88.120 ;
        RECT 101.640 87.835 101.980 88.085 ;
        RECT 102.150 87.525 102.320 88.755 ;
        RECT 102.820 88.545 103.030 89.400 ;
        RECT 101.640 87.275 102.320 87.525 ;
        RECT 100.865 86.855 101.970 87.105 ;
        RECT 97.810 86.450 100.125 86.535 ;
        RECT 93.140 85.970 93.840 86.180 ;
        RECT 89.985 84.920 91.095 85.360 ;
        RECT 91.265 85.090 91.800 85.345 ;
        RECT 89.985 84.730 91.460 84.920 ;
        RECT 89.985 84.715 90.590 84.730 ;
        RECT 87.220 84.170 88.415 84.420 ;
        RECT 88.735 84.365 90.590 84.715 ;
        RECT 91.270 84.590 91.460 84.730 ;
        RECT 91.630 84.805 91.800 85.090 ;
        RECT 91.980 84.975 92.460 85.360 ;
        RECT 92.655 84.805 92.920 85.340 ;
        RECT 91.630 84.550 92.920 84.805 ;
        RECT 86.880 83.740 87.505 84.000 ;
        RECT 86.880 83.565 87.050 83.740 ;
        RECT 84.980 83.520 85.880 83.555 ;
        RECT 77.930 82.770 80.800 83.520 ;
        RECT 80.970 83.000 83.720 83.520 ;
        RECT 83.890 83.300 85.880 83.520 ;
        RECT 80.970 82.770 83.180 83.000 ;
        RECT 83.890 82.830 85.150 83.300 ;
        RECT 86.065 83.130 87.050 83.565 ;
        RECT 87.700 83.560 88.415 84.170 ;
        RECT 87.220 83.300 88.415 83.560 ;
        RECT 85.325 82.870 87.505 83.130 ;
        RECT 85.325 82.840 87.050 82.870 ;
        RECT 75.530 82.310 76.990 82.770 ;
        RECT 74.100 82.140 75.360 82.200 ;
        RECT 73.300 81.740 73.890 81.990 ;
        RECT 74.100 81.570 75.880 82.140 ;
        RECT 73.300 81.390 75.880 81.570 ;
        RECT 76.050 81.390 76.990 82.310 ;
        RECT 79.540 82.600 80.800 82.770 ;
        RECT 79.540 81.850 81.320 82.600 ;
        RECT 81.490 82.310 83.180 82.770 ;
        RECT 83.350 82.670 85.150 82.830 ;
        RECT 83.350 82.400 85.895 82.670 ;
        RECT 86.065 82.400 87.050 82.840 ;
        RECT 87.700 82.775 88.415 83.300 ;
        RECT 89.985 83.890 90.590 84.365 ;
        RECT 90.760 84.075 91.100 84.550 ;
        RECT 91.630 84.365 91.800 84.550 ;
        RECT 91.335 84.115 91.800 84.365 ;
        RECT 89.985 83.675 91.435 83.890 ;
        RECT 91.630 83.785 91.800 84.115 ;
        RECT 91.980 84.150 92.920 84.380 ;
        RECT 93.140 84.155 93.310 85.970 ;
        RECT 94.220 85.695 94.550 86.400 ;
        RECT 94.755 85.865 95.130 86.420 ;
        RECT 95.860 86.190 96.030 86.450 ;
        RECT 95.360 85.875 96.030 86.190 ;
        RECT 95.860 85.810 96.030 85.875 ;
        RECT 98.580 86.195 100.125 86.450 ;
        RECT 100.865 86.265 101.470 86.855 ;
        RECT 102.140 86.685 102.320 87.275 ;
        RECT 101.640 86.435 102.320 86.685 ;
        RECT 93.590 85.525 95.560 85.695 ;
        RECT 93.590 84.910 93.760 85.525 ;
        RECT 93.930 85.035 95.220 85.355 ;
        RECT 93.930 84.890 94.260 85.035 ;
        RECT 93.590 84.505 93.760 84.740 ;
        RECT 94.470 84.675 95.190 84.865 ;
        RECT 95.390 84.810 95.560 85.525 ;
        RECT 95.860 85.520 97.000 85.810 ;
        RECT 98.580 85.640 99.295 86.195 ;
        RECT 95.860 84.950 96.030 85.520 ;
        RECT 96.200 85.140 98.030 85.350 ;
        RECT 98.200 85.310 99.295 85.640 ;
        RECT 96.200 85.120 98.410 85.140 ;
        RECT 97.840 84.950 98.410 85.120 ;
        RECT 95.860 84.620 96.445 84.950 ;
        RECT 96.745 84.780 97.670 84.950 ;
        RECT 98.580 84.780 99.295 85.310 ;
        RECT 95.360 84.505 95.690 84.585 ;
        RECT 93.590 84.335 95.690 84.505 ;
        RECT 91.980 83.970 92.475 84.150 ;
        RECT 93.140 83.970 93.810 84.155 ;
        RECT 92.645 83.785 93.810 83.970 ;
        RECT 93.990 83.875 94.290 84.335 ;
        RECT 95.860 84.165 96.030 84.620 ;
        RECT 96.745 84.610 98.010 84.780 ;
        RECT 96.745 84.430 96.975 84.610 ;
        RECT 94.470 83.995 94.800 84.165 ;
        RECT 95.060 83.995 96.030 84.165 ;
        RECT 96.200 84.115 96.975 84.430 ;
        RECT 97.255 84.115 97.670 84.440 ;
        RECT 97.840 84.230 98.010 84.610 ;
        RECT 98.220 84.450 99.295 84.780 ;
        RECT 100.865 86.015 101.970 86.265 ;
        RECT 100.865 85.160 101.470 86.015 ;
        RECT 102.140 85.845 102.320 86.435 ;
        RECT 102.490 88.375 103.030 88.545 ;
        RECT 103.200 89.055 103.850 89.420 ;
        RECT 104.020 89.180 104.570 89.510 ;
        RECT 104.740 89.275 106.070 89.505 ;
        RECT 103.200 88.545 103.380 89.055 ;
        RECT 104.020 88.885 104.190 89.180 ;
        RECT 104.740 89.010 104.910 89.275 ;
        RECT 103.550 88.715 104.190 88.885 ;
        RECT 104.450 88.840 104.910 89.010 ;
        RECT 105.080 88.755 105.730 89.105 ;
        RECT 105.900 89.010 106.070 89.275 ;
        RECT 106.240 89.320 106.910 89.510 ;
        RECT 108.220 89.420 108.550 89.540 ;
        RECT 106.240 89.180 107.630 89.320 ;
        RECT 105.900 88.840 106.570 89.010 ;
        RECT 106.740 88.990 107.630 89.180 ;
        RECT 107.800 89.250 108.830 89.420 ;
        RECT 109.000 89.410 109.290 89.710 ;
        RECT 109.460 89.755 110.175 90.130 ;
        RECT 109.460 89.415 111.005 89.755 ;
        RECT 104.020 88.580 104.190 88.715 ;
        RECT 106.740 88.580 106.910 88.990 ;
        RECT 107.800 88.780 107.970 89.250 ;
        RECT 102.490 86.405 102.660 88.375 ;
        RECT 103.200 88.215 103.850 88.545 ;
        RECT 102.830 86.700 103.030 88.150 ;
        RECT 104.020 88.045 105.480 88.580 ;
        RECT 103.200 87.875 105.480 88.045 ;
        RECT 104.020 87.830 105.480 87.875 ;
        RECT 105.650 88.310 106.910 88.580 ;
        RECT 107.250 88.480 107.970 88.780 ;
        RECT 108.220 88.750 108.470 89.080 ;
        RECT 105.650 88.030 107.580 88.310 ;
        RECT 108.220 88.145 108.470 88.520 ;
        RECT 103.200 87.235 103.850 87.565 ;
        RECT 103.200 86.725 103.380 87.235 ;
        RECT 104.020 87.065 104.960 87.830 ;
        RECT 105.650 87.660 106.910 88.030 ;
        RECT 107.780 87.830 108.470 88.145 ;
        RECT 108.640 88.360 108.830 89.250 ;
        RECT 109.460 89.240 110.175 89.415 ;
        RECT 109.000 88.990 110.175 89.240 ;
        RECT 108.640 88.030 109.190 88.360 ;
        RECT 103.550 86.910 104.960 87.065 ;
        RECT 105.130 86.910 106.910 87.660 ;
        RECT 103.550 86.895 104.190 86.910 ;
        RECT 103.200 86.475 103.850 86.725 ;
        RECT 102.490 86.235 103.030 86.405 ;
        RECT 102.820 85.930 103.030 86.235 ;
        RECT 101.640 85.760 102.320 85.845 ;
        RECT 103.210 85.760 103.460 86.305 ;
        RECT 101.640 85.530 103.460 85.760 ;
        RECT 103.630 85.550 103.850 86.475 ;
        RECT 104.020 86.310 104.190 86.895 ;
        RECT 106.740 86.740 106.910 86.910 ;
        RECT 109.460 86.740 110.175 88.990 ;
        RECT 111.745 87.935 112.350 91.340 ;
        RECT 110.495 87.585 112.350 87.935 ;
        RECT 104.450 86.480 104.910 86.650 ;
        RECT 104.020 85.980 104.570 86.310 ;
        RECT 104.740 86.215 104.910 86.480 ;
        RECT 105.080 86.385 105.730 86.735 ;
        RECT 105.900 86.480 106.570 86.650 ;
        RECT 106.740 86.480 107.920 86.740 ;
        RECT 105.900 86.215 106.070 86.480 ;
        RECT 106.740 86.310 106.910 86.480 ;
        RECT 108.100 86.310 108.620 86.740 ;
        RECT 108.800 86.465 110.175 86.740 ;
        RECT 104.740 85.985 106.070 86.215 ;
        RECT 106.240 85.980 106.910 86.310 ;
        RECT 107.080 86.295 108.620 86.310 ;
        RECT 107.080 86.140 109.290 86.295 ;
        RECT 107.080 86.035 107.750 86.140 ;
        RECT 108.100 86.125 109.290 86.140 ;
        RECT 108.830 86.045 109.290 86.125 ;
        RECT 104.020 85.370 104.190 85.980 ;
        RECT 106.740 85.835 106.910 85.980 ;
        RECT 109.460 85.995 110.175 86.465 ;
        RECT 111.745 85.995 112.350 87.585 ;
        RECT 104.450 85.625 106.570 85.810 ;
        RECT 106.740 85.620 107.755 85.835 ;
        RECT 107.950 85.725 108.550 85.955 ;
        RECT 109.460 85.870 109.630 85.995 ;
        RECT 108.965 85.820 109.630 85.870 ;
        RECT 112.180 85.820 112.350 85.995 ;
        RECT 100.865 84.880 102.140 85.160 ;
        RECT 102.340 85.045 103.030 85.360 ;
        RECT 100.865 84.715 101.470 84.880 ;
        RECT 97.840 84.040 98.410 84.230 ;
        RECT 89.985 83.030 90.590 83.675 ;
        RECT 91.630 83.555 92.230 83.785 ;
        RECT 92.645 83.640 93.310 83.785 ;
        RECT 93.990 83.675 94.320 83.875 ;
        RECT 94.540 83.825 94.800 83.995 ;
        RECT 90.760 83.370 91.430 83.475 ;
        RECT 92.510 83.385 92.970 83.465 ;
        RECT 91.780 83.370 92.970 83.385 ;
        RECT 90.760 83.215 92.970 83.370 ;
        RECT 90.760 83.200 92.300 83.215 ;
        RECT 89.985 82.775 91.600 83.030 ;
        RECT 87.700 82.700 87.870 82.775 ;
        RECT 87.220 82.400 87.870 82.700 ;
        RECT 83.350 82.310 85.150 82.400 ;
        RECT 81.490 82.140 82.430 82.310 ;
        RECT 81.490 81.850 82.910 82.140 ;
        RECT 79.540 81.680 79.710 81.850 ;
        RECT 73.300 81.320 74.270 81.390 ;
        RECT 72.540 80.940 73.130 81.110 ;
        RECT 73.300 80.980 73.930 81.150 ;
        RECT 74.100 81.115 74.270 81.320 ;
        RECT 73.300 80.730 73.470 80.980 ;
        RECT 74.100 80.945 74.730 81.115 ;
        RECT 74.100 80.770 74.270 80.945 ;
        RECT 74.900 80.790 76.250 81.220 ;
        RECT 76.820 81.195 76.990 81.390 ;
        RECT 76.420 80.865 76.990 81.195 ;
        RECT 77.210 81.125 77.475 81.660 ;
        RECT 77.670 81.295 78.150 81.680 ;
        RECT 78.330 81.410 78.865 81.665 ;
        RECT 78.330 81.125 78.500 81.410 ;
        RECT 79.035 81.240 79.710 81.680 ;
        RECT 77.210 80.870 78.500 81.125 ;
        RECT 78.670 81.220 79.710 81.240 ;
        RECT 82.260 81.810 82.910 81.850 ;
        RECT 83.095 81.815 83.670 82.130 ;
        RECT 84.980 82.120 85.150 82.310 ;
        RECT 87.700 82.130 87.870 82.400 ;
        RECT 84.015 81.860 84.810 82.080 ;
        RECT 78.670 81.050 80.215 81.220 ;
        RECT 78.670 80.910 78.860 81.050 ;
        RECT 74.900 80.775 75.070 80.790 ;
        RECT 71.380 80.475 72.010 80.730 ;
        RECT 72.180 80.475 73.470 80.730 ;
        RECT 73.640 80.520 74.270 80.770 ;
        RECT 65.480 80.060 67.400 80.300 ;
        RECT 62.750 80.030 63.390 80.060 ;
        RECT 60.840 79.720 61.360 79.780 ;
        RECT 62.165 79.720 62.950 79.850 ;
        RECT 60.840 79.545 62.950 79.720 ;
        RECT 63.220 79.360 63.390 80.030 ;
        RECT 63.985 79.890 65.350 79.945 ;
        RECT 63.560 79.775 65.660 79.890 ;
        RECT 63.560 79.640 64.115 79.775 ;
        RECT 65.220 79.720 65.660 79.775 ;
        RECT 60.500 79.090 61.305 79.360 ;
        RECT 62.265 79.090 63.390 79.360 ;
        RECT 60.500 78.920 60.670 79.090 ;
        RECT 63.220 78.920 63.390 79.090 ;
        RECT 60.500 78.630 61.395 78.920 ;
        RECT 62.055 78.630 63.390 78.920 ;
        RECT 60.500 78.460 60.670 78.630 ;
        RECT 63.220 78.460 63.390 78.630 ;
        RECT 60.500 76.875 61.215 78.460 ;
        RECT 62.785 78.155 63.390 78.460 ;
        RECT 63.665 78.495 63.835 79.430 ;
        RECT 64.305 79.365 64.900 79.605 ;
        RECT 65.490 79.555 65.660 79.720 ;
        RECT 65.940 79.780 67.400 80.060 ;
        RECT 67.570 80.210 68.830 80.300 ;
        RECT 67.570 79.895 69.330 80.210 ;
        RECT 65.070 79.195 65.290 79.550 ;
        RECT 64.005 79.025 65.290 79.195 ;
        RECT 64.005 78.665 64.370 79.025 ;
        RECT 65.490 78.855 65.660 79.360 ;
        RECT 64.540 78.685 65.660 78.855 ;
        RECT 65.940 79.090 66.860 79.780 ;
        RECT 67.570 79.610 68.830 79.895 ;
        RECT 69.560 79.885 69.935 80.440 ;
        RECT 70.140 79.715 70.470 80.420 ;
        RECT 71.380 80.260 71.550 80.475 ;
        RECT 71.380 80.200 72.370 80.260 ;
        RECT 70.850 80.030 72.370 80.200 ;
        RECT 70.850 79.990 71.550 80.030 ;
        RECT 67.030 79.090 68.830 79.610 ;
        RECT 65.940 78.920 66.110 79.090 ;
        RECT 68.660 78.920 68.830 79.090 ;
        RECT 64.540 78.495 64.710 78.685 ;
        RECT 63.665 78.325 64.710 78.495 ;
        RECT 65.940 78.630 66.835 78.920 ;
        RECT 67.495 78.630 68.830 78.920 ;
        RECT 69.130 79.545 71.100 79.715 ;
        RECT 69.130 78.830 69.300 79.545 ;
        RECT 69.470 79.055 70.760 79.375 ;
        RECT 70.430 78.910 70.760 79.055 ;
        RECT 70.930 78.930 71.100 79.545 ;
        RECT 71.380 79.360 71.550 79.990 ;
        RECT 72.540 79.950 72.790 80.280 ;
        RECT 74.100 80.275 74.270 80.520 ;
        RECT 74.440 80.445 75.070 80.775 ;
        RECT 76.080 80.695 76.250 80.790 ;
        RECT 75.240 80.450 75.910 80.620 ;
        RECT 76.080 80.525 76.520 80.695 ;
        RECT 74.100 80.260 75.070 80.275 ;
        RECT 72.960 80.105 75.070 80.260 ;
        RECT 72.960 80.030 74.270 80.105 ;
        RECT 71.720 79.780 72.350 79.860 ;
        RECT 72.950 79.780 73.930 79.860 ;
        RECT 71.720 79.530 73.930 79.780 ;
        RECT 74.100 79.360 74.270 80.030 ;
        RECT 75.240 79.700 75.410 80.450 ;
        RECT 76.820 80.355 76.990 80.865 ;
        RECT 77.210 80.470 78.150 80.700 ;
        RECT 76.310 80.290 76.990 80.355 ;
        RECT 77.655 80.290 78.150 80.470 ;
        RECT 78.330 80.685 78.500 80.870 ;
        RECT 78.330 80.435 78.795 80.685 ;
        RECT 75.580 79.870 76.140 80.280 ;
        RECT 76.310 80.040 77.485 80.290 ;
        RECT 78.330 80.105 78.500 80.435 ;
        RECT 79.030 80.395 79.370 80.870 ;
        RECT 79.540 80.780 80.215 81.050 ;
        RECT 80.385 80.950 80.920 81.205 ;
        RECT 79.540 80.590 80.580 80.780 ;
        RECT 79.540 80.210 79.710 80.590 ;
        RECT 80.390 80.450 80.580 80.590 ;
        RECT 80.750 80.665 80.920 80.950 ;
        RECT 81.100 80.835 81.580 81.220 ;
        RECT 81.775 80.665 82.040 81.200 ;
        RECT 80.750 80.410 82.040 80.665 ;
        RECT 82.260 80.460 82.430 81.810 ;
        RECT 82.710 81.245 83.670 81.625 ;
        RECT 84.015 81.190 84.280 81.860 ;
        RECT 84.980 81.790 85.950 82.120 ;
        RECT 86.975 81.800 87.870 82.130 ;
        RECT 84.980 81.690 85.150 81.790 ;
        RECT 84.470 81.360 85.150 81.690 ;
        RECT 87.190 81.615 87.360 81.620 ;
        RECT 84.015 80.965 84.810 81.190 ;
        RECT 84.980 81.110 85.150 81.360 ;
        RECT 85.320 81.610 87.445 81.615 ;
        RECT 85.320 81.440 87.490 81.610 ;
        RECT 85.320 81.280 86.290 81.440 ;
        RECT 86.980 81.280 87.490 81.440 ;
        RECT 82.600 80.680 83.170 80.870 ;
        RECT 76.820 79.960 77.485 80.040 ;
        RECT 76.310 79.700 76.650 79.810 ;
        RECT 75.240 79.520 76.650 79.700 ;
        RECT 71.380 79.150 72.370 79.360 ;
        RECT 72.960 79.150 74.270 79.360 ;
        RECT 75.065 79.160 75.410 79.520 ;
        RECT 76.820 79.365 76.990 79.960 ;
        RECT 77.900 79.875 78.500 80.105 ;
        RECT 78.695 79.995 79.710 80.210 ;
        RECT 77.160 79.705 77.620 79.785 ;
        RECT 77.160 79.690 78.350 79.705 ;
        RECT 78.700 79.690 79.370 79.795 ;
        RECT 77.160 79.535 79.370 79.690 ;
        RECT 77.830 79.520 79.370 79.535 ;
        RECT 79.540 79.750 79.710 79.995 ;
        RECT 79.880 79.935 80.220 80.410 ;
        RECT 80.750 80.225 80.920 80.410 ;
        RECT 80.455 79.975 80.920 80.225 ;
        RECT 79.540 79.535 80.555 79.750 ;
        RECT 80.750 79.645 80.920 79.975 ;
        RECT 81.100 80.010 82.040 80.240 ;
        RECT 82.260 80.130 82.790 80.460 ;
        RECT 83.000 80.300 83.170 80.680 ;
        RECT 83.340 80.470 83.755 80.795 ;
        RECT 84.035 80.480 84.810 80.795 ;
        RECT 84.980 80.780 85.950 81.110 ;
        RECT 86.470 81.100 86.710 81.270 ;
        RECT 87.700 81.110 87.870 81.800 ;
        RECT 90.420 82.770 91.600 82.775 ;
        RECT 91.780 82.770 92.300 83.200 ;
        RECT 93.140 83.045 93.310 83.640 ;
        RECT 94.540 83.655 95.585 83.825 ;
        RECT 94.540 83.465 94.710 83.655 ;
        RECT 92.480 82.770 93.310 83.045 ;
        RECT 93.590 83.295 94.710 83.465 ;
        RECT 93.590 82.790 93.760 83.295 ;
        RECT 94.880 83.125 95.245 83.485 ;
        RECT 93.960 82.955 95.245 83.125 ;
        RECT 90.420 82.600 90.590 82.770 ;
        RECT 90.420 82.160 91.095 82.600 ;
        RECT 91.265 82.330 91.800 82.585 ;
        RECT 90.420 81.970 91.460 82.160 ;
        RECT 90.420 81.680 90.590 81.970 ;
        RECT 91.270 81.830 91.460 81.970 ;
        RECT 91.630 82.045 91.800 82.330 ;
        RECT 91.980 82.215 92.460 82.600 ;
        RECT 92.655 82.045 92.920 82.580 ;
        RECT 91.630 81.790 92.920 82.045 ;
        RECT 93.140 82.090 93.310 82.770 ;
        RECT 93.960 82.600 94.180 82.955 ;
        RECT 93.590 82.430 93.760 82.595 ;
        RECT 94.350 82.545 94.945 82.785 ;
        RECT 95.415 82.720 95.585 83.655 ;
        RECT 95.860 83.550 96.030 83.995 ;
        RECT 96.200 83.720 96.995 83.945 ;
        RECT 95.860 83.220 96.540 83.550 ;
        RECT 95.860 82.540 96.030 83.220 ;
        RECT 96.730 83.050 96.995 83.720 ;
        RECT 97.340 83.285 98.300 83.665 ;
        RECT 98.580 83.100 99.295 84.450 ;
        RECT 99.615 84.365 101.470 84.715 ;
        RECT 101.810 84.410 102.530 84.710 ;
        RECT 102.780 84.670 103.030 85.045 ;
        RECT 103.200 84.830 103.750 85.160 ;
        RECT 104.020 85.120 104.650 85.370 ;
        RECT 104.820 85.175 105.770 85.455 ;
        RECT 106.740 85.385 106.910 85.620 ;
        RECT 106.280 85.120 106.910 85.385 ;
        RECT 96.200 82.830 96.995 83.050 ;
        RECT 97.340 82.780 97.915 83.095 ;
        RECT 98.100 82.775 99.295 83.100 ;
        RECT 100.865 84.200 101.470 84.365 ;
        RECT 100.865 83.870 102.190 84.200 ;
        RECT 102.360 83.940 102.530 84.410 ;
        RECT 102.780 84.110 103.030 84.440 ;
        RECT 103.200 83.940 103.390 84.830 ;
        RECT 104.020 84.200 104.190 85.120 ;
        RECT 104.780 84.950 106.145 85.005 ;
        RECT 104.470 84.835 106.570 84.950 ;
        RECT 104.470 84.780 104.910 84.835 ;
        RECT 104.470 84.615 104.640 84.780 ;
        RECT 106.015 84.700 106.570 84.835 ;
        RECT 106.740 84.780 106.910 85.120 ;
        RECT 107.080 84.960 107.420 85.435 ;
        RECT 107.950 85.395 108.120 85.725 ;
        RECT 108.965 85.540 110.175 85.820 ;
        RECT 107.655 85.145 108.120 85.395 ;
        RECT 107.950 84.960 108.120 85.145 ;
        RECT 108.300 85.360 108.795 85.540 ;
        RECT 108.300 85.130 109.240 85.360 ;
        RECT 107.590 84.780 107.780 84.920 ;
        RECT 103.560 83.950 104.190 84.200 ;
        RECT 100.865 83.060 101.470 83.870 ;
        RECT 102.360 83.770 103.390 83.940 ;
        RECT 101.640 83.480 102.190 83.680 ;
        RECT 102.780 83.650 103.110 83.770 ;
        RECT 103.560 83.480 103.850 83.780 ;
        RECT 101.640 83.230 103.850 83.480 ;
        RECT 104.020 83.425 104.190 83.950 ;
        RECT 104.470 83.915 104.640 84.420 ;
        RECT 104.840 84.255 105.060 84.610 ;
        RECT 105.230 84.425 105.825 84.665 ;
        RECT 106.740 84.590 107.780 84.780 ;
        RECT 107.950 84.705 109.240 84.960 ;
        RECT 104.840 84.085 106.125 84.255 ;
        RECT 104.470 83.745 105.590 83.915 ;
        RECT 105.420 83.555 105.590 83.745 ;
        RECT 105.760 83.725 106.125 84.085 ;
        RECT 106.295 83.555 106.465 84.490 ;
        RECT 104.020 83.060 104.690 83.425 ;
        RECT 100.865 82.775 102.610 83.060 ;
        RECT 98.100 82.770 98.750 82.775 ;
        RECT 98.580 82.540 98.750 82.770 ;
        RECT 93.590 82.375 94.030 82.430 ;
        RECT 95.135 82.375 95.690 82.510 ;
        RECT 93.590 82.260 95.690 82.375 ;
        RECT 95.860 82.330 97.170 82.540 ;
        RECT 97.760 82.330 98.750 82.540 ;
        RECT 93.900 82.205 95.265 82.260 ;
        RECT 95.860 82.090 96.030 82.330 ;
        RECT 93.140 81.840 93.770 82.090 ;
        RECT 86.120 80.875 86.710 81.100 ;
        RECT 86.895 80.875 87.870 81.110 ;
        RECT 84.035 80.300 84.265 80.480 ;
        RECT 83.000 80.130 84.265 80.300 ;
        RECT 84.980 80.290 85.150 80.780 ;
        RECT 86.120 80.380 86.290 80.875 ;
        RECT 86.460 80.445 87.370 80.705 ;
        RECT 81.100 79.830 81.595 80.010 ;
        RECT 82.260 79.830 82.430 80.130 ;
        RECT 83.340 79.960 84.265 80.130 ;
        RECT 84.565 79.960 85.150 80.290 ;
        RECT 85.320 80.130 86.290 80.380 ;
        RECT 87.700 80.290 87.870 80.875 ;
        RECT 88.090 81.125 88.355 81.660 ;
        RECT 88.550 81.295 89.030 81.680 ;
        RECT 89.210 81.410 89.745 81.665 ;
        RECT 89.210 81.125 89.380 81.410 ;
        RECT 89.915 81.240 90.590 81.680 ;
        RECT 90.760 81.315 91.100 81.790 ;
        RECT 91.630 81.605 91.800 81.790 ;
        RECT 91.335 81.355 91.800 81.605 ;
        RECT 88.090 80.870 89.380 81.125 ;
        RECT 89.550 81.130 90.590 81.240 ;
        RECT 89.550 81.050 91.435 81.130 ;
        RECT 89.550 80.910 89.740 81.050 ;
        RECT 90.420 80.915 91.435 81.050 ;
        RECT 91.630 81.025 91.800 81.355 ;
        RECT 91.980 81.390 92.920 81.620 ;
        RECT 91.980 81.210 92.475 81.390 ;
        RECT 93.140 81.230 93.310 81.840 ;
        RECT 93.940 81.755 94.890 82.035 ;
        RECT 95.400 81.825 96.030 82.090 ;
        RECT 96.200 81.910 98.410 82.160 ;
        RECT 96.200 81.830 97.180 81.910 ;
        RECT 97.780 81.830 98.410 81.910 ;
        RECT 98.580 82.140 98.750 82.330 ;
        RECT 101.300 82.770 102.610 82.775 ;
        RECT 103.220 83.055 104.690 83.060 ;
        RECT 104.870 83.335 105.200 83.535 ;
        RECT 105.420 83.385 106.465 83.555 ;
        RECT 106.740 84.150 107.415 84.590 ;
        RECT 107.950 84.420 108.120 84.705 ;
        RECT 107.585 84.165 108.120 84.420 ;
        RECT 108.300 84.150 108.780 84.535 ;
        RECT 108.975 84.170 109.240 84.705 ;
        RECT 109.460 84.235 110.175 85.540 ;
        RECT 106.740 83.875 106.910 84.150 ;
        RECT 106.740 83.705 107.370 83.875 ;
        RECT 103.220 82.770 104.190 83.055 ;
        RECT 104.870 82.875 105.170 83.335 ;
        RECT 105.420 83.215 105.680 83.385 ;
        RECT 106.740 83.215 106.910 83.705 ;
        RECT 107.540 83.550 108.890 83.980 ;
        RECT 109.460 83.955 111.005 84.235 ;
        RECT 109.060 83.895 111.005 83.955 ;
        RECT 109.060 83.625 110.175 83.895 ;
        RECT 107.540 83.535 107.710 83.550 ;
        RECT 105.350 83.045 105.680 83.215 ;
        RECT 105.940 83.045 106.910 83.215 ;
        RECT 107.080 83.205 107.710 83.535 ;
        RECT 108.720 83.455 108.890 83.550 ;
        RECT 107.880 83.210 108.550 83.380 ;
        RECT 108.720 83.285 109.160 83.455 ;
        RECT 106.740 83.035 106.910 83.045 ;
        RECT 101.300 82.140 101.470 82.770 ;
        RECT 98.580 81.865 99.410 82.140 ;
        RECT 95.860 81.660 96.030 81.825 ;
        RECT 93.570 81.400 95.690 81.585 ;
        RECT 95.860 81.430 97.170 81.660 ;
        RECT 95.860 81.230 96.030 81.430 ;
        RECT 97.340 81.410 97.590 81.740 ;
        RECT 98.580 81.660 98.750 81.865 ;
        RECT 99.590 81.710 100.110 82.140 ;
        RECT 100.290 81.880 101.470 82.140 ;
        RECT 101.640 81.880 102.310 82.050 ;
        RECT 101.300 81.710 101.470 81.880 ;
        RECT 99.590 81.695 101.130 81.710 ;
        RECT 97.760 81.430 98.750 81.660 ;
        RECT 98.920 81.540 101.130 81.695 ;
        RECT 98.920 81.525 100.110 81.540 ;
        RECT 98.920 81.445 99.380 81.525 ;
        RECT 100.460 81.435 101.130 81.540 ;
        RECT 93.140 81.210 93.690 81.230 ;
        RECT 88.090 80.470 89.030 80.700 ;
        RECT 88.535 80.290 89.030 80.470 ;
        RECT 89.210 80.685 89.380 80.870 ;
        RECT 89.210 80.435 89.675 80.685 ;
        RECT 86.480 80.135 87.370 80.265 ;
        RECT 76.820 79.350 77.650 79.365 ;
        RECT 75.580 79.155 76.140 79.350 ;
        RECT 75.630 79.150 75.800 79.155 ;
        RECT 71.380 78.920 71.550 79.150 ;
        RECT 74.100 78.920 74.270 79.150 ;
        RECT 76.310 79.110 77.650 79.350 ;
        RECT 76.820 79.090 77.650 79.110 ;
        RECT 77.830 79.090 78.350 79.520 ;
        RECT 79.540 79.350 79.710 79.535 ;
        RECT 80.750 79.415 81.350 79.645 ;
        RECT 81.765 79.600 82.430 79.830 ;
        RECT 82.600 79.790 83.170 79.960 ;
        RECT 84.980 79.945 85.150 79.960 ;
        RECT 82.600 79.770 84.810 79.790 ;
        RECT 81.765 79.500 82.810 79.600 ;
        RECT 82.980 79.560 84.810 79.770 ;
        RECT 84.980 79.615 85.870 79.945 ;
        RECT 78.530 79.090 79.710 79.350 ;
        RECT 76.820 78.920 76.990 79.090 ;
        RECT 79.540 78.920 79.710 79.090 ;
        RECT 79.880 79.230 80.550 79.335 ;
        RECT 81.630 79.245 82.090 79.325 ;
        RECT 80.900 79.230 82.090 79.245 ;
        RECT 79.880 79.075 82.090 79.230 ;
        RECT 82.260 79.270 82.810 79.500 ;
        RECT 84.980 79.390 85.150 79.615 ;
        RECT 86.120 79.395 86.290 80.130 ;
        RECT 86.460 79.965 87.370 80.135 ;
        RECT 87.700 79.960 88.365 80.290 ;
        RECT 89.210 80.105 89.380 80.435 ;
        RECT 89.910 80.395 90.250 80.870 ;
        RECT 90.420 80.270 90.590 80.915 ;
        RECT 91.630 80.795 92.230 81.025 ;
        RECT 92.645 80.900 93.690 81.210 ;
        RECT 93.860 80.995 95.190 81.225 ;
        RECT 92.645 80.880 93.310 80.900 ;
        RECT 90.760 80.610 91.430 80.715 ;
        RECT 92.510 80.625 92.970 80.705 ;
        RECT 91.780 80.610 92.970 80.625 ;
        RECT 90.760 80.455 92.970 80.610 ;
        RECT 90.760 80.440 92.300 80.455 ;
        RECT 90.420 80.210 91.600 80.270 ;
        RECT 86.460 79.435 87.365 79.790 ;
        RECT 79.880 79.060 81.420 79.075 ;
        RECT 69.500 78.695 70.220 78.885 ;
        RECT 64.450 78.155 64.710 78.325 ;
        RECT 64.930 78.275 65.260 78.475 ;
        RECT 65.940 78.460 66.110 78.630 ;
        RECT 68.660 78.460 68.830 78.630 ;
        RECT 65.940 78.365 66.655 78.460 ;
        RECT 62.785 77.985 64.190 78.155 ;
        RECT 64.450 77.985 64.780 78.155 ;
        RECT 60.500 76.535 62.045 76.875 ;
        RECT 60.500 73.115 61.215 76.535 ;
        RECT 62.785 76.275 63.390 77.985 ;
        RECT 64.960 77.815 65.260 78.275 ;
        RECT 65.440 77.995 66.655 78.365 ;
        RECT 63.560 77.645 65.660 77.815 ;
        RECT 63.560 77.565 63.890 77.645 ;
        RECT 63.690 76.625 63.860 77.340 ;
        RECT 64.060 77.285 64.780 77.475 ;
        RECT 65.490 77.410 65.660 77.645 ;
        RECT 64.990 77.115 65.320 77.260 ;
        RECT 64.030 76.795 65.320 77.115 ;
        RECT 65.490 76.625 65.660 77.240 ;
        RECT 63.690 76.455 65.660 76.625 ;
        RECT 65.940 76.875 66.655 77.995 ;
        RECT 68.225 78.185 68.830 78.460 ;
        RECT 69.000 78.525 69.330 78.605 ;
        RECT 70.930 78.525 71.100 78.760 ;
        RECT 69.000 78.355 71.100 78.525 ;
        RECT 71.380 78.630 72.275 78.920 ;
        RECT 72.935 78.630 74.705 78.920 ;
        RECT 71.380 78.460 71.550 78.630 ;
        RECT 74.100 78.460 74.705 78.630 ;
        RECT 68.225 78.015 69.630 78.185 ;
        RECT 69.890 78.015 70.220 78.185 ;
        RECT 65.940 76.535 67.485 76.875 ;
        RECT 62.785 75.960 63.890 76.275 ;
        RECT 62.785 75.220 63.390 75.960 ;
        RECT 64.120 75.730 64.495 76.285 ;
        RECT 64.700 75.750 65.030 76.455 ;
        RECT 65.940 76.180 66.655 76.535 ;
        RECT 65.410 75.970 66.655 76.180 ;
        RECT 63.560 75.580 64.495 75.730 ;
        RECT 65.200 75.580 65.725 75.710 ;
        RECT 63.560 75.390 65.725 75.580 ;
        RECT 64.700 75.380 65.725 75.390 ;
        RECT 62.785 75.055 64.400 75.220 ;
        RECT 61.535 75.050 64.400 75.055 ;
        RECT 61.535 74.705 63.390 75.050 ;
        RECT 62.785 74.380 63.390 74.705 ;
        RECT 63.605 74.705 64.530 74.880 ;
        RECT 64.700 74.830 65.030 75.380 ;
        RECT 65.940 75.210 66.655 75.970 ;
        RECT 65.330 75.040 66.655 75.210 ;
        RECT 68.225 76.110 68.830 78.015 ;
        RECT 69.890 77.845 70.150 78.015 ;
        RECT 70.400 77.895 70.700 78.355 ;
        RECT 71.380 78.175 72.095 78.460 ;
        RECT 69.105 77.675 70.150 77.845 ;
        RECT 70.370 77.695 70.700 77.895 ;
        RECT 70.880 77.805 72.095 78.175 ;
        RECT 69.105 76.740 69.275 77.675 ;
        RECT 69.445 77.145 69.810 77.505 ;
        RECT 69.980 77.485 70.150 77.675 ;
        RECT 69.980 77.315 71.100 77.485 ;
        RECT 69.445 76.975 70.730 77.145 ;
        RECT 69.745 76.565 70.340 76.805 ;
        RECT 70.510 76.620 70.730 76.975 ;
        RECT 70.930 76.810 71.100 77.315 ;
        RECT 71.380 76.875 72.095 77.805 ;
        RECT 69.000 76.395 69.555 76.530 ;
        RECT 70.930 76.450 71.100 76.615 ;
        RECT 70.660 76.395 71.100 76.450 ;
        RECT 69.000 76.280 71.100 76.395 ;
        RECT 71.380 76.535 72.925 76.875 ;
        RECT 69.425 76.225 70.790 76.280 ;
        RECT 71.380 76.110 72.095 76.535 ;
        RECT 68.225 75.845 69.290 76.110 ;
        RECT 68.225 75.250 68.830 75.845 ;
        RECT 69.800 75.775 70.750 76.055 ;
        RECT 70.920 75.860 72.095 76.110 ;
        RECT 69.000 75.420 71.120 75.605 ;
        RECT 71.380 75.250 72.095 75.860 ;
        RECT 68.225 75.055 69.330 75.250 ;
        RECT 65.200 74.715 65.720 74.870 ;
        RECT 63.605 74.660 64.580 74.705 ;
        RECT 65.160 74.660 65.720 74.715 ;
        RECT 63.605 74.550 65.720 74.660 ;
        RECT 64.450 74.540 65.720 74.550 ;
        RECT 64.450 74.490 65.285 74.540 ;
        RECT 62.785 74.210 64.305 74.380 ;
        RECT 65.940 74.370 66.655 75.040 ;
        RECT 66.975 74.920 69.330 75.055 ;
        RECT 69.500 75.015 70.830 75.245 ;
        RECT 66.975 74.705 68.830 74.920 ;
        RECT 69.500 74.750 69.670 75.015 ;
        RECT 62.785 73.860 63.390 74.210 ;
        RECT 65.425 74.200 66.655 74.370 ;
        RECT 65.940 73.860 66.655 74.200 ;
        RECT 62.785 73.115 63.825 73.860 ;
        RECT 60.500 72.940 60.670 73.115 ;
        RECT 63.220 72.940 63.825 73.115 ;
        RECT 60.500 71.355 61.215 72.940 ;
        RECT 60.500 71.015 62.045 71.355 ;
        RECT 60.500 67.595 61.215 71.015 ;
        RECT 62.785 70.455 63.825 72.940 ;
        RECT 65.395 73.115 66.655 73.860 ;
        RECT 68.225 74.320 68.830 74.705 ;
        RECT 69.000 74.580 69.670 74.750 ;
        RECT 69.840 74.495 70.490 74.845 ;
        RECT 70.660 74.750 70.830 75.015 ;
        RECT 71.000 74.920 72.095 75.250 ;
        RECT 73.665 75.515 74.705 78.460 ;
        RECT 76.275 78.630 77.715 78.920 ;
        RECT 78.375 78.890 79.710 78.920 ;
        RECT 78.375 78.630 80.720 78.890 ;
        RECT 80.900 78.630 81.420 79.060 ;
        RECT 82.260 78.920 82.430 79.270 ;
        RECT 84.010 79.100 85.150 79.390 ;
        RECT 85.320 79.215 86.290 79.395 ;
        RECT 87.700 79.365 87.870 79.960 ;
        RECT 88.780 79.875 89.380 80.105 ;
        RECT 89.575 80.010 91.600 80.210 ;
        RECT 91.780 80.010 92.300 80.440 ;
        RECT 93.140 80.300 93.310 80.880 ;
        RECT 93.860 80.730 94.030 80.995 ;
        RECT 93.570 80.560 94.030 80.730 ;
        RECT 94.200 80.475 94.850 80.825 ;
        RECT 95.020 80.730 95.190 80.995 ;
        RECT 95.360 81.220 96.030 81.230 ;
        RECT 98.580 81.270 98.750 81.430 ;
        RECT 101.300 81.380 101.970 81.710 ;
        RECT 102.140 81.615 102.310 81.880 ;
        RECT 102.480 81.785 103.130 82.135 ;
        RECT 103.300 81.880 103.760 82.050 ;
        RECT 103.300 81.615 103.470 81.880 ;
        RECT 104.020 81.710 104.190 82.770 ;
        RECT 104.470 82.705 106.570 82.875 ;
        RECT 104.470 82.470 104.640 82.705 ;
        RECT 106.240 82.625 106.570 82.705 ;
        RECT 106.740 82.865 107.710 83.035 ;
        RECT 105.350 82.345 106.070 82.535 ;
        RECT 102.140 81.385 103.470 81.615 ;
        RECT 103.640 81.380 104.190 81.710 ;
        RECT 104.470 81.685 104.640 82.300 ;
        RECT 104.810 82.175 105.140 82.320 ;
        RECT 104.810 81.855 106.100 82.175 ;
        RECT 106.270 81.685 106.440 82.400 ;
        RECT 104.470 81.515 106.440 81.685 ;
        RECT 106.740 81.680 106.910 82.865 ;
        RECT 107.880 82.460 108.050 83.210 ;
        RECT 109.460 83.115 110.175 83.625 ;
        RECT 108.220 82.630 108.780 83.040 ;
        RECT 108.950 82.800 110.175 83.115 ;
        RECT 108.950 82.460 109.290 82.570 ;
        RECT 107.880 82.280 109.290 82.460 ;
        RECT 107.705 81.920 108.050 82.280 ;
        RECT 109.460 82.110 110.175 82.800 ;
        RECT 111.745 82.415 112.350 85.820 ;
        RECT 108.220 81.915 108.780 82.110 ;
        RECT 108.270 81.910 108.440 81.915 ;
        RECT 108.950 81.870 110.175 82.110 ;
        RECT 110.495 82.065 112.350 82.415 ;
        RECT 109.460 81.680 110.175 81.870 ;
        RECT 98.580 81.220 99.245 81.270 ;
        RECT 95.360 80.900 97.120 81.220 ;
        RECT 95.020 80.560 95.690 80.730 ;
        RECT 95.860 80.300 97.120 80.900 ;
        RECT 97.290 80.940 99.245 81.220 ;
        RECT 99.660 81.125 100.260 81.355 ;
        RECT 101.300 81.235 101.470 81.380 ;
        RECT 97.290 80.470 98.750 80.940 ;
        RECT 99.415 80.760 99.910 80.940 ;
        RECT 98.970 80.530 99.910 80.760 ;
        RECT 100.090 80.795 100.260 81.125 ;
        RECT 100.455 81.020 101.470 81.235 ;
        RECT 104.020 81.240 104.190 81.380 ;
        RECT 101.640 81.025 103.760 81.210 ;
        RECT 104.020 81.030 104.720 81.240 ;
        RECT 100.090 80.545 100.555 80.795 ;
        RECT 93.140 80.285 94.600 80.300 ;
        RECT 92.480 80.010 94.600 80.285 ;
        RECT 89.575 79.995 90.590 80.010 ;
        RECT 88.040 79.705 88.500 79.785 ;
        RECT 88.040 79.690 89.230 79.705 ;
        RECT 89.580 79.690 90.250 79.795 ;
        RECT 88.040 79.535 90.250 79.690 ;
        RECT 88.710 79.520 90.250 79.535 ;
        RECT 85.320 79.145 87.530 79.215 ;
        RECT 84.980 78.970 85.150 79.100 ;
        RECT 86.120 79.045 87.530 79.145 ;
        RECT 84.980 78.920 85.530 78.970 ;
        RECT 82.260 78.905 83.155 78.920 ;
        RECT 81.600 78.630 83.155 78.905 ;
        RECT 83.815 78.640 85.530 78.920 ;
        RECT 85.710 78.670 87.030 78.875 ;
        RECT 87.200 78.720 87.530 79.045 ;
        RECT 87.700 79.090 88.530 79.365 ;
        RECT 88.710 79.090 89.230 79.520 ;
        RECT 90.420 79.380 90.590 79.995 ;
        RECT 93.140 79.780 94.600 80.010 ;
        RECT 90.420 79.350 91.095 79.380 ;
        RECT 89.410 79.090 91.095 79.350 ;
        RECT 91.265 79.110 91.800 79.365 ;
        RECT 87.700 78.920 87.870 79.090 ;
        RECT 90.420 78.940 91.095 79.090 ;
        RECT 90.420 78.920 91.460 78.940 ;
        RECT 83.815 78.630 85.150 78.640 ;
        RECT 76.275 78.030 76.990 78.630 ;
        RECT 79.540 78.460 79.710 78.630 ;
        RECT 77.250 78.200 77.710 78.370 ;
        RECT 76.275 77.700 77.370 78.030 ;
        RECT 77.540 77.935 77.710 78.200 ;
        RECT 77.880 78.105 78.530 78.455 ;
        RECT 78.700 78.200 79.370 78.370 ;
        RECT 79.540 78.200 80.850 78.460 ;
        RECT 78.700 77.935 78.870 78.200 ;
        RECT 79.540 78.030 79.710 78.200 ;
        RECT 77.540 77.705 78.870 77.935 ;
        RECT 79.040 77.700 79.710 78.030 ;
        RECT 79.880 77.700 80.850 78.030 ;
        RECT 81.020 77.700 81.270 78.460 ;
        RECT 81.460 78.120 82.090 78.460 ;
        RECT 76.275 77.335 76.990 77.700 ;
        RECT 79.540 77.530 79.710 77.700 ;
        RECT 77.250 77.345 79.370 77.530 ;
        RECT 79.540 77.360 80.510 77.530 ;
        RECT 75.445 77.090 76.990 77.335 ;
        RECT 75.445 76.995 77.450 77.090 ;
        RECT 76.275 76.840 77.450 76.995 ;
        RECT 77.620 76.895 78.570 77.175 ;
        RECT 79.540 77.105 79.710 77.360 ;
        RECT 80.680 77.190 80.850 77.700 ;
        RECT 81.460 77.610 81.630 78.120 ;
        RECT 82.260 77.950 82.430 78.630 ;
        RECT 84.980 78.460 85.150 78.630 ;
        RECT 87.700 78.630 88.595 78.920 ;
        RECT 89.255 78.750 91.460 78.920 ;
        RECT 89.255 78.630 90.590 78.750 ;
        RECT 84.980 78.020 85.655 78.460 ;
        RECT 85.825 78.190 86.360 78.445 ;
        RECT 81.800 77.780 82.430 77.950 ;
        RECT 79.080 76.840 79.710 77.105 ;
        RECT 79.880 76.860 80.850 77.190 ;
        RECT 73.665 75.165 75.955 75.515 ;
        RECT 73.665 75.055 74.705 75.165 ;
        RECT 70.660 74.580 71.120 74.750 ;
        RECT 68.225 73.880 69.335 74.320 ;
        RECT 69.505 74.050 70.040 74.305 ;
        RECT 68.225 73.690 69.700 73.880 ;
        RECT 68.225 73.115 68.830 73.690 ;
        RECT 69.510 73.550 69.700 73.690 ;
        RECT 69.870 73.765 70.040 74.050 ;
        RECT 70.220 73.935 70.700 74.320 ;
        RECT 70.895 73.765 71.160 74.300 ;
        RECT 69.870 73.510 71.160 73.765 ;
        RECT 65.395 72.940 66.110 73.115 ;
        RECT 68.660 72.940 68.830 73.115 ;
        RECT 69.000 73.035 69.340 73.510 ;
        RECT 69.870 73.325 70.040 73.510 ;
        RECT 69.575 73.075 70.040 73.325 ;
        RECT 65.395 72.275 66.655 72.940 ;
        RECT 64.565 71.935 66.655 72.275 ;
        RECT 65.395 71.355 66.655 71.935 ;
        RECT 68.225 72.850 68.830 72.940 ;
        RECT 68.225 72.635 69.675 72.850 ;
        RECT 69.870 72.745 70.040 73.075 ;
        RECT 70.220 73.110 71.160 73.340 ;
        RECT 71.380 73.115 72.095 74.920 ;
        RECT 72.415 74.705 74.705 75.055 ;
        RECT 73.665 73.575 74.705 74.705 ;
        RECT 76.275 75.145 76.990 76.840 ;
        RECT 77.580 76.670 78.945 76.725 ;
        RECT 79.540 76.690 79.710 76.840 ;
        RECT 77.270 76.555 79.370 76.670 ;
        RECT 77.270 76.500 77.710 76.555 ;
        RECT 77.270 76.335 77.440 76.500 ;
        RECT 78.815 76.420 79.370 76.555 ;
        RECT 79.540 76.435 80.510 76.690 ;
        RECT 80.680 76.610 80.850 76.860 ;
        RECT 81.020 76.780 81.270 77.530 ;
        RECT 81.460 77.360 82.090 77.610 ;
        RECT 81.440 76.610 81.690 77.190 ;
        RECT 81.880 76.770 82.090 77.360 ;
        RECT 77.270 75.635 77.440 76.140 ;
        RECT 77.640 75.975 77.860 76.330 ;
        RECT 78.030 76.145 78.625 76.385 ;
        RECT 77.640 75.805 78.925 75.975 ;
        RECT 77.270 75.465 78.390 75.635 ;
        RECT 78.220 75.275 78.390 75.465 ;
        RECT 78.560 75.445 78.925 75.805 ;
        RECT 79.095 75.275 79.265 76.210 ;
        RECT 76.275 74.775 77.490 75.145 ;
        RECT 77.670 75.055 78.000 75.255 ;
        RECT 78.220 75.105 79.265 75.275 ;
        RECT 79.540 76.160 79.710 76.435 ;
        RECT 80.680 76.330 81.690 76.610 ;
        RECT 81.860 76.440 82.090 76.770 ;
        RECT 82.260 77.570 82.430 77.780 ;
        RECT 82.690 77.740 83.150 77.910 ;
        RECT 82.260 77.240 82.810 77.570 ;
        RECT 82.980 77.475 83.150 77.740 ;
        RECT 83.320 77.645 83.970 77.995 ;
        RECT 84.140 77.740 84.810 77.910 ;
        RECT 84.980 77.830 86.020 78.020 ;
        RECT 84.140 77.475 84.310 77.740 ;
        RECT 84.980 77.570 85.150 77.830 ;
        RECT 85.830 77.690 86.020 77.830 ;
        RECT 86.190 77.905 86.360 78.190 ;
        RECT 86.540 78.075 87.020 78.460 ;
        RECT 87.215 77.905 87.480 78.440 ;
        RECT 86.190 77.650 87.480 77.905 ;
        RECT 87.700 78.400 87.870 78.630 ;
        RECT 90.420 78.400 90.590 78.630 ;
        RECT 91.270 78.610 91.460 78.750 ;
        RECT 91.630 78.825 91.800 79.110 ;
        RECT 91.980 78.995 92.460 79.380 ;
        RECT 92.655 78.825 92.920 79.360 ;
        RECT 91.630 78.570 92.920 78.825 ;
        RECT 93.140 79.090 94.060 79.780 ;
        RECT 94.770 79.610 97.640 80.300 ;
        RECT 94.230 79.550 97.640 79.610 ;
        RECT 97.810 79.550 98.750 80.470 ;
        RECT 100.090 80.360 100.260 80.545 ;
        RECT 100.790 80.360 101.130 80.835 ;
        RECT 101.300 80.785 101.470 81.020 ;
        RECT 101.300 80.520 101.930 80.785 ;
        RECT 102.440 80.575 103.390 80.855 ;
        RECT 104.020 80.770 104.190 81.030 ;
        RECT 105.100 80.810 105.430 81.515 ;
        RECT 105.635 80.790 106.010 81.345 ;
        RECT 106.740 81.335 107.345 81.680 ;
        RECT 106.240 81.020 107.345 81.335 ;
        RECT 103.560 80.520 104.190 80.770 ;
        RECT 98.970 80.105 100.260 80.360 ;
        RECT 98.970 79.570 99.235 80.105 ;
        RECT 99.430 79.550 99.910 79.935 ;
        RECT 100.090 79.820 100.260 80.105 ;
        RECT 100.430 80.180 100.620 80.320 ;
        RECT 101.300 80.180 101.470 80.520 ;
        RECT 102.065 80.350 103.430 80.405 ;
        RECT 100.430 79.990 101.470 80.180 ;
        RECT 101.640 80.235 103.740 80.350 ;
        RECT 101.640 80.100 102.195 80.235 ;
        RECT 103.300 80.180 103.740 80.235 ;
        RECT 100.090 79.565 100.625 79.820 ;
        RECT 100.795 79.550 101.470 79.990 ;
        RECT 94.230 79.275 96.030 79.550 ;
        RECT 94.230 79.090 96.830 79.275 ;
        RECT 93.140 78.920 93.310 79.090 ;
        RECT 95.860 79.020 96.830 79.090 ;
        RECT 97.000 79.100 98.010 79.380 ;
        RECT 95.860 78.920 96.030 79.020 ;
        RECT 93.140 78.630 94.035 78.920 ;
        RECT 94.695 78.630 96.030 78.920 ;
        RECT 97.000 78.850 97.170 79.100 ;
        RECT 87.700 78.190 88.690 78.400 ;
        RECT 89.280 78.190 90.590 78.400 ;
        RECT 82.980 77.245 84.310 77.475 ;
        RECT 84.480 77.240 85.150 77.570 ;
        RECT 82.260 76.630 82.430 77.240 ;
        RECT 82.690 76.885 84.810 77.070 ;
        RECT 84.980 76.990 85.150 77.240 ;
        RECT 85.320 77.175 85.660 77.650 ;
        RECT 86.190 77.465 86.360 77.650 ;
        RECT 87.700 77.520 87.870 78.190 ;
        RECT 88.040 77.770 90.250 78.020 ;
        RECT 88.040 77.690 88.670 77.770 ;
        RECT 89.270 77.690 90.250 77.770 ;
        RECT 90.420 77.910 90.590 78.190 ;
        RECT 90.760 78.095 91.100 78.570 ;
        RECT 91.630 78.385 91.800 78.570 ;
        RECT 91.335 78.135 91.800 78.385 ;
        RECT 90.420 77.695 91.435 77.910 ;
        RECT 91.630 77.805 91.800 78.135 ;
        RECT 91.980 78.170 92.920 78.400 ;
        RECT 91.980 77.990 92.475 78.170 ;
        RECT 93.140 77.990 93.310 78.630 ;
        RECT 95.860 78.350 96.030 78.630 ;
        RECT 96.200 78.520 97.170 78.850 ;
        RECT 95.860 78.180 96.830 78.350 ;
        RECT 85.895 77.215 86.360 77.465 ;
        RECT 84.980 76.775 85.995 76.990 ;
        RECT 86.190 76.885 86.360 77.215 ;
        RECT 86.540 77.250 87.480 77.480 ;
        RECT 87.700 77.290 88.690 77.520 ;
        RECT 86.540 77.070 87.035 77.250 ;
        RECT 87.700 77.070 87.870 77.290 ;
        RECT 88.860 77.270 89.110 77.600 ;
        RECT 90.420 77.520 90.590 77.695 ;
        RECT 91.630 77.575 92.230 77.805 ;
        RECT 92.645 77.660 93.310 77.990 ;
        RECT 93.570 77.740 94.030 77.910 ;
        RECT 89.280 77.290 90.590 77.520 ;
        RECT 93.140 77.570 93.310 77.660 ;
        RECT 82.260 76.380 82.890 76.630 ;
        RECT 83.060 76.435 84.010 76.715 ;
        RECT 84.980 76.645 85.150 76.775 ;
        RECT 86.190 76.655 86.790 76.885 ;
        RECT 87.205 76.740 87.870 77.070 ;
        RECT 88.130 76.820 88.590 76.990 ;
        RECT 84.520 76.380 85.150 76.645 ;
        RECT 87.700 76.650 87.870 76.740 ;
        RECT 82.260 76.160 82.430 76.380 ;
        RECT 83.020 76.210 84.385 76.265 ;
        RECT 76.275 73.575 76.990 74.775 ;
        RECT 77.670 74.595 77.970 75.055 ;
        RECT 78.220 74.935 78.480 75.105 ;
        RECT 79.540 74.935 80.145 76.160 ;
        RECT 78.150 74.765 78.480 74.935 ;
        RECT 78.740 74.765 80.145 74.935 ;
        RECT 77.270 74.425 79.370 74.595 ;
        RECT 77.270 74.190 77.440 74.425 ;
        RECT 79.040 74.345 79.370 74.425 ;
        RECT 78.150 74.065 78.870 74.255 ;
        RECT 73.665 73.400 74.270 73.575 ;
        RECT 76.820 73.400 76.990 73.575 ;
        RECT 73.665 73.115 74.705 73.400 ;
        RECT 70.220 72.930 70.715 73.110 ;
        RECT 71.380 72.940 71.550 73.115 ;
        RECT 74.100 72.940 74.705 73.115 ;
        RECT 71.380 72.930 72.095 72.940 ;
        RECT 68.225 71.990 68.830 72.635 ;
        RECT 69.870 72.515 70.470 72.745 ;
        RECT 70.885 72.600 72.095 72.930 ;
        RECT 69.000 72.420 69.670 72.435 ;
        RECT 69.000 72.330 69.680 72.420 ;
        RECT 70.750 72.345 71.210 72.425 ;
        RECT 70.020 72.330 71.210 72.345 ;
        RECT 69.000 72.175 71.210 72.330 ;
        RECT 69.000 72.160 70.540 72.175 ;
        RECT 68.225 71.730 69.840 71.990 ;
        RECT 70.020 71.730 70.540 72.160 ;
        RECT 71.380 72.005 72.095 72.600 ;
        RECT 70.720 71.730 72.095 72.005 ;
        RECT 68.225 71.560 68.830 71.730 ;
        RECT 71.380 71.560 72.095 71.730 ;
        RECT 65.395 71.015 67.485 71.355 ;
        RECT 62.785 70.105 65.075 70.455 ;
        RECT 62.785 69.535 63.825 70.105 ;
        RECT 61.535 69.185 63.825 69.535 ;
        RECT 62.785 68.515 63.825 69.185 ;
        RECT 65.395 68.515 66.655 71.015 ;
        RECT 68.225 69.740 69.920 71.560 ;
        RECT 70.090 71.355 72.095 71.560 ;
        RECT 70.090 71.015 72.925 71.355 ;
        RECT 70.090 69.910 72.095 71.015 ;
        RECT 68.225 69.535 70.440 69.740 ;
        RECT 66.975 69.185 70.440 69.535 ;
        RECT 62.785 68.340 63.390 68.515 ;
        RECT 65.940 68.340 66.655 68.515 ;
        RECT 62.785 67.650 64.480 68.340 ;
        RECT 64.650 67.820 66.655 68.340 ;
        RECT 62.785 67.595 65.020 67.650 ;
        RECT 60.500 66.960 60.670 67.595 ;
        RECT 63.220 67.130 65.020 67.595 ;
        RECT 65.190 67.595 66.655 67.820 ;
        RECT 68.225 68.050 70.440 69.185 ;
        RECT 70.610 68.050 72.095 69.910 ;
        RECT 73.665 69.995 74.705 72.940 ;
        RECT 76.275 72.960 76.990 73.400 ;
        RECT 77.270 73.405 77.440 74.020 ;
        RECT 77.610 73.895 77.940 74.040 ;
        RECT 77.610 73.575 78.900 73.895 ;
        RECT 79.070 73.405 79.240 74.120 ;
        RECT 77.270 73.235 79.240 73.405 ;
        RECT 76.275 72.750 77.520 72.960 ;
        RECT 76.275 71.990 76.990 72.750 ;
        RECT 77.900 72.530 78.230 73.235 ;
        RECT 78.435 72.510 78.810 73.065 ;
        RECT 79.540 73.055 80.145 74.765 ;
        RECT 81.715 74.685 82.430 76.160 ;
        RECT 82.710 76.095 84.810 76.210 ;
        RECT 82.710 76.040 83.150 76.095 ;
        RECT 82.710 75.875 82.880 76.040 ;
        RECT 84.255 75.960 84.810 76.095 ;
        RECT 84.980 76.130 85.150 76.380 ;
        RECT 85.320 76.470 85.990 76.575 ;
        RECT 87.070 76.485 87.530 76.565 ;
        RECT 86.340 76.470 87.530 76.485 ;
        RECT 85.320 76.315 87.530 76.470 ;
        RECT 87.700 76.320 88.250 76.650 ;
        RECT 88.420 76.555 88.590 76.820 ;
        RECT 88.760 76.725 89.410 77.075 ;
        RECT 90.420 77.050 90.590 77.290 ;
        RECT 90.760 77.390 91.430 77.495 ;
        RECT 92.510 77.405 92.970 77.485 ;
        RECT 91.780 77.390 92.970 77.405 ;
        RECT 90.760 77.235 92.970 77.390 ;
        RECT 93.140 77.240 93.690 77.570 ;
        RECT 93.860 77.475 94.030 77.740 ;
        RECT 94.200 77.645 94.850 77.995 ;
        RECT 95.020 77.740 95.690 77.910 ;
        RECT 95.020 77.475 95.190 77.740 ;
        RECT 95.860 77.570 96.030 78.180 ;
        RECT 97.000 78.010 97.170 78.520 ;
        RECT 97.340 78.180 97.590 78.930 ;
        RECT 97.760 78.520 98.010 79.100 ;
        RECT 98.180 78.940 98.410 79.270 ;
        RECT 98.200 78.350 98.410 78.940 ;
        RECT 97.780 78.100 98.410 78.350 ;
        RECT 98.580 78.920 98.750 79.550 ;
        RECT 101.300 78.920 101.470 79.550 ;
        RECT 98.580 78.630 99.475 78.920 ;
        RECT 100.135 78.630 101.470 78.920 ;
        RECT 101.745 78.955 101.915 79.890 ;
        RECT 102.385 79.825 102.980 80.065 ;
        RECT 103.570 80.015 103.740 80.180 ;
        RECT 104.020 80.270 104.190 80.520 ;
        RECT 104.405 80.640 104.930 80.770 ;
        RECT 105.635 80.640 106.570 80.790 ;
        RECT 104.405 80.450 106.570 80.640 ;
        RECT 104.405 80.440 105.430 80.450 ;
        RECT 104.020 80.100 104.800 80.270 ;
        RECT 103.150 79.655 103.370 80.010 ;
        RECT 102.085 79.485 103.370 79.655 ;
        RECT 102.085 79.125 102.450 79.485 ;
        RECT 103.570 79.315 103.740 79.820 ;
        RECT 102.620 79.145 103.740 79.315 ;
        RECT 104.020 79.430 104.190 80.100 ;
        RECT 104.410 79.775 104.930 79.930 ;
        RECT 105.100 79.890 105.430 80.440 ;
        RECT 106.740 80.280 107.345 81.020 ;
        RECT 105.730 80.110 107.345 80.280 ;
        RECT 104.410 79.720 104.970 79.775 ;
        RECT 105.600 79.765 106.525 79.940 ;
        RECT 105.550 79.720 106.525 79.765 ;
        RECT 104.410 79.610 106.525 79.720 ;
        RECT 104.410 79.600 105.680 79.610 ;
        RECT 104.845 79.550 105.680 79.600 ;
        RECT 106.740 79.440 107.345 80.110 ;
        RECT 108.915 80.475 110.175 81.680 ;
        RECT 111.745 80.475 112.350 82.065 ;
        RECT 108.915 80.300 109.630 80.475 ;
        RECT 112.180 80.300 112.350 80.475 ;
        RECT 108.915 80.095 110.920 80.300 ;
        RECT 108.085 79.780 110.920 80.095 ;
        RECT 108.085 79.755 110.380 79.780 ;
        RECT 104.020 79.260 104.705 79.430 ;
        RECT 105.825 79.270 107.345 79.440 ;
        RECT 102.620 78.955 102.790 79.145 ;
        RECT 101.745 78.785 102.790 78.955 ;
        RECT 98.580 78.435 98.750 78.630 ;
        RECT 101.300 78.615 101.470 78.630 ;
        RECT 102.530 78.615 102.790 78.785 ;
        RECT 103.010 78.735 103.340 78.935 ;
        RECT 104.020 78.920 104.190 79.260 ;
        RECT 106.740 78.920 107.345 79.270 ;
        RECT 104.020 78.825 104.915 78.920 ;
        RECT 98.580 78.105 99.150 78.435 ;
        RECT 96.200 77.680 97.170 78.010 ;
        RECT 93.860 77.245 95.190 77.475 ;
        RECT 95.360 77.510 96.030 77.570 ;
        RECT 95.360 77.250 97.170 77.510 ;
        RECT 97.340 77.250 97.590 78.010 ;
        RECT 97.780 77.590 97.950 78.100 ;
        RECT 98.580 77.930 98.750 78.105 ;
        RECT 99.320 78.030 100.670 78.460 ;
        RECT 101.300 78.445 102.270 78.615 ;
        RECT 102.530 78.445 102.860 78.615 ;
        RECT 101.300 78.355 101.470 78.445 ;
        RECT 100.840 78.185 101.470 78.355 ;
        RECT 103.040 78.275 103.340 78.735 ;
        RECT 103.520 78.630 104.915 78.825 ;
        RECT 105.575 78.630 107.345 78.920 ;
        RECT 103.520 78.455 104.190 78.630 ;
        RECT 106.740 78.460 107.345 78.630 ;
        RECT 99.320 77.935 99.490 78.030 ;
        RECT 98.120 77.760 98.750 77.930 ;
        RECT 99.050 77.765 99.490 77.935 ;
        RECT 100.500 78.015 100.670 78.030 ;
        RECT 98.580 77.595 98.750 77.760 ;
        RECT 99.660 77.690 100.330 77.860 ;
        RECT 97.780 77.250 98.410 77.590 ;
        RECT 98.580 77.280 99.260 77.595 ;
        RECT 95.360 77.240 96.030 77.250 ;
        RECT 90.760 77.220 92.300 77.235 ;
        RECT 89.580 76.820 90.250 76.990 ;
        RECT 89.580 76.555 89.750 76.820 ;
        RECT 90.420 76.790 91.600 77.050 ;
        RECT 91.780 76.790 92.300 77.220 ;
        RECT 93.140 77.065 93.310 77.240 ;
        RECT 92.480 76.790 93.310 77.065 ;
        RECT 93.570 76.885 95.690 77.070 ;
        RECT 90.420 76.650 90.590 76.790 ;
        RECT 88.420 76.325 89.750 76.555 ;
        RECT 89.920 76.620 90.590 76.650 ;
        RECT 93.140 76.630 93.310 76.790 ;
        RECT 93.140 76.620 93.770 76.630 ;
        RECT 89.920 76.320 91.025 76.620 ;
        RECT 85.320 76.300 86.860 76.315 ;
        RECT 82.710 75.175 82.880 75.680 ;
        RECT 83.080 75.515 83.300 75.870 ;
        RECT 83.470 75.685 84.065 75.925 ;
        RECT 84.980 75.870 86.160 76.130 ;
        RECT 86.340 75.870 86.860 76.300 ;
        RECT 87.700 76.145 87.870 76.320 ;
        RECT 87.040 75.870 87.870 76.145 ;
        RECT 88.130 75.965 90.250 76.150 ;
        RECT 83.080 75.345 84.365 75.515 ;
        RECT 82.710 75.005 83.830 75.175 ;
        RECT 83.660 74.815 83.830 75.005 ;
        RECT 84.000 74.985 84.365 75.345 ;
        RECT 84.535 74.815 84.705 75.750 ;
        RECT 81.715 74.575 82.930 74.685 ;
        RECT 80.885 74.315 82.930 74.575 ;
        RECT 83.110 74.595 83.440 74.795 ;
        RECT 83.660 74.645 84.705 74.815 ;
        RECT 84.980 75.595 85.150 75.870 ;
        RECT 87.700 75.710 87.870 75.870 ;
        RECT 84.980 75.425 85.610 75.595 ;
        RECT 84.980 74.755 85.150 75.425 ;
        RECT 85.780 75.270 87.130 75.700 ;
        RECT 87.700 75.675 88.330 75.710 ;
        RECT 87.300 75.460 88.330 75.675 ;
        RECT 88.500 75.515 89.450 75.795 ;
        RECT 90.420 75.725 91.025 76.320 ;
        RECT 89.960 75.460 91.025 75.725 ;
        RECT 87.300 75.345 87.870 75.460 ;
        RECT 85.780 75.255 85.950 75.270 ;
        RECT 85.320 74.925 85.950 75.255 ;
        RECT 86.960 75.175 87.130 75.270 ;
        RECT 86.120 74.930 86.790 75.100 ;
        RECT 86.960 75.005 87.400 75.175 ;
        RECT 80.885 74.235 82.430 74.315 ;
        RECT 79.040 72.755 80.145 73.055 ;
        RECT 79.040 72.740 81.395 72.755 ;
        RECT 77.205 72.360 77.730 72.490 ;
        RECT 78.435 72.360 79.370 72.510 ;
        RECT 77.205 72.170 79.370 72.360 ;
        RECT 79.540 72.405 81.395 72.740 ;
        RECT 81.715 72.500 82.430 74.235 ;
        RECT 83.110 74.135 83.410 74.595 ;
        RECT 83.660 74.475 83.920 74.645 ;
        RECT 84.980 74.585 85.950 74.755 ;
        RECT 84.980 74.475 85.150 74.585 ;
        RECT 83.590 74.305 83.920 74.475 ;
        RECT 84.180 74.305 85.150 74.475 ;
        RECT 82.710 73.965 84.810 74.135 ;
        RECT 82.710 73.730 82.880 73.965 ;
        RECT 84.480 73.885 84.810 73.965 ;
        RECT 83.590 73.605 84.310 73.795 ;
        RECT 82.710 72.945 82.880 73.560 ;
        RECT 83.050 73.435 83.380 73.580 ;
        RECT 83.050 73.115 84.340 73.435 ;
        RECT 84.510 72.945 84.680 73.660 ;
        RECT 82.710 72.775 84.680 72.945 ;
        RECT 84.980 73.360 85.150 74.305 ;
        RECT 86.120 74.180 86.290 74.930 ;
        RECT 87.700 74.835 87.870 75.345 ;
        RECT 88.460 75.290 89.825 75.345 ;
        RECT 88.150 75.175 90.250 75.290 ;
        RECT 88.150 75.120 88.590 75.175 ;
        RECT 88.150 74.955 88.320 75.120 ;
        RECT 89.695 75.040 90.250 75.175 ;
        RECT 86.460 74.350 87.020 74.760 ;
        RECT 87.190 74.520 87.870 74.835 ;
        RECT 87.190 74.180 87.530 74.290 ;
        RECT 86.120 74.000 87.530 74.180 ;
        RECT 85.945 73.640 86.290 74.000 ;
        RECT 87.700 73.830 87.870 74.520 ;
        RECT 88.150 74.255 88.320 74.760 ;
        RECT 88.520 74.595 88.740 74.950 ;
        RECT 88.910 74.765 89.505 75.005 ;
        RECT 88.520 74.425 89.805 74.595 ;
        RECT 88.150 74.085 89.270 74.255 ;
        RECT 89.100 73.895 89.270 74.085 ;
        RECT 89.440 74.065 89.805 74.425 ;
        RECT 89.975 73.895 90.145 74.830 ;
        RECT 86.460 73.635 87.020 73.830 ;
        RECT 87.190 73.765 87.870 73.830 ;
        RECT 86.510 73.630 86.680 73.635 ;
        RECT 87.190 73.590 88.370 73.765 ;
        RECT 87.700 73.395 88.370 73.590 ;
        RECT 88.550 73.675 88.880 73.875 ;
        RECT 89.100 73.725 90.145 73.895 ;
        RECT 84.980 73.130 86.290 73.360 ;
        RECT 77.205 72.160 78.230 72.170 ;
        RECT 76.275 71.820 77.600 71.990 ;
        RECT 76.275 71.815 76.990 71.820 ;
        RECT 75.445 71.475 76.990 71.815 ;
        RECT 76.275 71.150 76.990 71.475 ;
        RECT 77.210 71.495 77.730 71.650 ;
        RECT 77.900 71.610 78.230 72.160 ;
        RECT 79.540 72.000 80.145 72.405 ;
        RECT 78.530 71.830 80.145 72.000 ;
        RECT 77.210 71.440 77.770 71.495 ;
        RECT 78.400 71.485 79.325 71.660 ;
        RECT 78.350 71.440 79.325 71.485 ;
        RECT 77.210 71.330 79.325 71.440 ;
        RECT 77.210 71.320 78.480 71.330 ;
        RECT 77.645 71.270 78.480 71.320 ;
        RECT 79.540 71.160 80.145 71.830 ;
        RECT 76.275 70.980 77.505 71.150 ;
        RECT 78.625 70.990 80.145 71.160 ;
        RECT 76.275 70.640 76.990 70.980 ;
        RECT 79.540 70.815 80.145 70.990 ;
        RECT 81.715 72.290 82.960 72.500 ;
        RECT 81.715 71.530 82.430 72.290 ;
        RECT 83.340 72.070 83.670 72.775 ;
        RECT 83.875 72.050 84.250 72.605 ;
        RECT 84.980 72.595 85.150 73.130 ;
        RECT 86.460 73.050 86.710 73.380 ;
        RECT 87.700 73.360 87.870 73.395 ;
        RECT 86.880 73.130 87.870 73.360 ;
        RECT 88.550 73.215 88.850 73.675 ;
        RECT 89.100 73.555 89.360 73.725 ;
        RECT 90.420 73.555 91.025 75.460 ;
        RECT 92.595 76.380 93.770 76.620 ;
        RECT 93.940 76.435 94.890 76.715 ;
        RECT 95.860 76.645 96.030 77.240 ;
        RECT 98.580 77.060 98.750 77.280 ;
        RECT 99.430 77.110 99.990 77.520 ;
        RECT 97.390 77.015 97.560 77.020 ;
        RECT 96.825 76.650 97.170 77.010 ;
        RECT 97.340 76.820 97.900 77.015 ;
        RECT 98.070 76.820 98.750 77.060 ;
        RECT 95.400 76.380 96.030 76.645 ;
        RECT 92.595 75.035 93.310 76.380 ;
        RECT 93.900 76.210 95.265 76.265 ;
        RECT 93.590 76.095 95.690 76.210 ;
        RECT 93.590 76.040 94.030 76.095 ;
        RECT 93.590 75.875 93.760 76.040 ;
        RECT 95.135 75.960 95.690 76.095 ;
        RECT 95.860 76.065 96.030 76.380 ;
        RECT 97.000 76.470 98.410 76.650 ;
        RECT 91.765 74.695 93.310 75.035 ;
        RECT 93.590 75.175 93.760 75.680 ;
        RECT 93.960 75.515 94.180 75.870 ;
        RECT 94.350 75.685 94.945 75.925 ;
        RECT 95.860 75.895 96.830 76.065 ;
        RECT 93.960 75.345 95.245 75.515 ;
        RECT 93.590 75.005 94.710 75.175 ;
        RECT 94.540 74.815 94.710 75.005 ;
        RECT 94.880 74.985 95.245 75.345 ;
        RECT 95.415 74.815 95.585 75.750 ;
        RECT 89.030 73.385 89.360 73.555 ;
        RECT 89.620 73.385 91.025 73.555 ;
        RECT 90.420 73.215 91.025 73.385 ;
        RECT 92.595 74.685 93.310 74.695 ;
        RECT 92.595 74.315 93.810 74.685 ;
        RECT 93.990 74.595 94.320 74.795 ;
        RECT 94.540 74.645 95.585 74.815 ;
        RECT 95.860 75.225 96.030 75.895 ;
        RECT 96.200 75.395 96.830 75.725 ;
        RECT 97.000 75.720 97.170 76.470 ;
        RECT 98.070 76.360 98.410 76.470 ;
        RECT 98.580 76.590 98.750 76.820 ;
        RECT 98.920 76.940 99.260 77.050 ;
        RECT 100.160 76.940 100.330 77.690 ;
        RECT 100.500 77.685 101.130 78.015 ;
        RECT 101.300 77.515 101.470 78.185 ;
        RECT 101.640 78.105 103.740 78.275 ;
        RECT 101.640 78.025 101.970 78.105 ;
        RECT 100.500 77.345 101.470 77.515 ;
        RECT 98.920 76.760 100.330 76.940 ;
        RECT 98.580 76.350 99.260 76.590 ;
        RECT 99.430 76.395 99.990 76.590 ;
        RECT 100.160 76.400 100.505 76.760 ;
        RECT 101.300 76.735 101.470 77.345 ;
        RECT 101.770 77.085 101.940 77.800 ;
        RECT 102.140 77.745 102.860 77.935 ;
        RECT 103.570 77.870 103.740 78.105 ;
        RECT 104.020 77.950 104.190 78.455 ;
        RECT 104.360 78.120 104.990 78.460 ;
        RECT 104.020 77.780 104.650 77.950 ;
        RECT 103.070 77.575 103.400 77.720 ;
        RECT 102.110 77.255 103.400 77.575 ;
        RECT 103.570 77.085 103.740 77.700 ;
        RECT 101.770 76.915 103.740 77.085 ;
        RECT 101.300 76.420 101.970 76.735 ;
        RECT 99.770 76.390 99.940 76.395 ;
        RECT 97.340 75.890 97.900 76.300 ;
        RECT 98.580 76.160 98.750 76.350 ;
        RECT 101.300 76.160 101.470 76.420 ;
        RECT 102.200 76.190 102.575 76.745 ;
        RECT 102.780 76.210 103.110 76.915 ;
        RECT 104.020 76.640 104.190 77.780 ;
        RECT 104.820 77.610 104.990 78.120 ;
        RECT 105.180 77.700 105.430 78.460 ;
        RECT 105.600 78.275 107.345 78.460 ;
        RECT 108.915 79.090 110.380 79.755 ;
        RECT 111.090 79.610 112.350 80.300 ;
        RECT 110.550 79.090 112.350 79.610 ;
        RECT 108.915 78.920 109.630 79.090 ;
        RECT 112.180 78.920 112.350 79.090 ;
        RECT 108.915 78.630 110.355 78.920 ;
        RECT 111.015 78.630 112.350 78.920 ;
        RECT 108.915 78.460 109.630 78.630 ;
        RECT 112.180 78.460 112.350 78.630 ;
        RECT 105.600 78.200 108.595 78.275 ;
        RECT 105.600 77.700 106.570 78.030 ;
        RECT 106.740 77.925 108.595 78.200 ;
        RECT 103.490 76.430 104.190 76.640 ;
        RECT 104.360 77.360 104.990 77.610 ;
        RECT 104.360 76.770 104.570 77.360 ;
        RECT 104.360 76.440 104.590 76.770 ;
        RECT 104.760 76.610 105.010 77.190 ;
        RECT 105.180 76.780 105.430 77.530 ;
        RECT 105.600 77.190 105.770 77.700 ;
        RECT 106.740 77.530 107.345 77.925 ;
        RECT 105.940 77.360 107.345 77.530 ;
        RECT 105.600 76.860 106.570 77.190 ;
        RECT 105.600 76.610 105.770 76.860 ;
        RECT 106.740 76.690 107.345 77.360 ;
        RECT 98.580 76.130 99.295 76.160 ;
        RECT 98.070 75.815 99.295 76.130 ;
        RECT 97.000 75.550 97.670 75.720 ;
        RECT 96.660 75.380 96.830 75.395 ;
        RECT 97.840 75.475 98.280 75.645 ;
        RECT 97.840 75.380 98.010 75.475 ;
        RECT 95.860 75.055 96.490 75.225 ;
        RECT 95.860 74.780 96.030 75.055 ;
        RECT 96.660 74.950 98.010 75.380 ;
        RECT 98.580 75.305 99.295 75.815 ;
        RECT 98.180 74.975 99.295 75.305 ;
        RECT 98.580 74.780 99.295 74.975 ;
        RECT 85.320 72.880 86.300 72.960 ;
        RECT 86.900 72.880 87.530 72.960 ;
        RECT 85.320 72.630 87.530 72.880 ;
        RECT 84.480 72.460 85.150 72.595 ;
        RECT 87.700 72.460 87.870 73.130 ;
        RECT 88.150 73.045 90.250 73.215 ;
        RECT 88.150 72.810 88.320 73.045 ;
        RECT 89.920 72.965 90.250 73.045 ;
        RECT 89.030 72.685 89.750 72.875 ;
        RECT 90.420 72.865 92.275 73.215 ;
        RECT 84.480 72.280 86.290 72.460 ;
        RECT 84.980 72.250 86.290 72.280 ;
        RECT 86.880 72.250 87.870 72.460 ;
        RECT 82.645 71.900 83.170 72.030 ;
        RECT 83.875 71.900 84.810 72.050 ;
        RECT 82.645 71.710 84.810 71.900 ;
        RECT 84.980 72.020 85.150 72.250 ;
        RECT 87.700 72.020 87.870 72.250 ;
        RECT 82.645 71.700 83.670 71.710 ;
        RECT 81.715 71.360 83.040 71.530 ;
        RECT 81.715 70.815 82.430 71.360 ;
        RECT 82.650 71.035 83.170 71.190 ;
        RECT 83.340 71.150 83.670 71.700 ;
        RECT 84.980 71.540 86.240 72.020 ;
        RECT 83.970 71.370 86.240 71.540 ;
        RECT 82.650 70.980 83.210 71.035 ;
        RECT 83.840 71.025 84.765 71.200 ;
        RECT 83.790 70.980 84.765 71.025 ;
        RECT 82.650 70.870 84.765 70.980 ;
        RECT 82.650 70.860 83.920 70.870 ;
        RECT 79.540 70.640 79.710 70.815 ;
        RECT 82.260 70.690 82.430 70.815 ;
        RECT 83.085 70.810 83.920 70.860 ;
        RECT 84.980 70.700 86.240 71.370 ;
        RECT 82.260 70.640 82.945 70.690 ;
        RECT 73.665 69.645 75.955 69.995 ;
        RECT 73.665 69.535 74.705 69.645 ;
        RECT 72.415 69.185 74.705 69.535 ;
        RECT 68.225 67.595 68.830 68.050 ;
        RECT 65.190 67.130 66.110 67.595 ;
        RECT 63.220 66.960 63.390 67.130 ;
        RECT 65.940 66.960 66.110 67.130 ;
        RECT 68.660 66.960 68.830 67.595 ;
        RECT 71.380 67.595 72.095 68.050 ;
        RECT 73.665 68.055 74.705 69.185 ;
        RECT 76.275 68.990 78.280 70.640 ;
        RECT 76.275 68.055 77.760 68.990 ;
        RECT 78.450 68.820 80.800 70.640 ;
        RECT 80.970 70.520 82.945 70.640 ;
        RECT 84.065 70.530 86.240 70.700 ;
        RECT 80.970 70.180 82.430 70.520 ;
        RECT 84.980 70.200 86.240 70.530 ;
        RECT 86.410 71.580 87.870 72.020 ;
        RECT 88.150 72.025 88.320 72.640 ;
        RECT 88.490 72.515 88.820 72.660 ;
        RECT 88.490 72.195 89.780 72.515 ;
        RECT 89.950 72.025 90.120 72.740 ;
        RECT 88.150 71.855 90.120 72.025 ;
        RECT 86.410 71.370 88.400 71.580 ;
        RECT 86.410 70.610 87.870 71.370 ;
        RECT 88.780 71.150 89.110 71.855 ;
        RECT 89.315 71.130 89.690 71.685 ;
        RECT 90.420 71.675 91.025 72.865 ;
        RECT 89.920 71.360 91.025 71.675 ;
        RECT 90.420 71.275 91.025 71.360 ;
        RECT 92.595 72.500 93.310 74.315 ;
        RECT 93.990 74.135 94.290 74.595 ;
        RECT 94.540 74.475 94.800 74.645 ;
        RECT 95.860 74.475 96.465 74.780 ;
        RECT 94.470 74.305 94.800 74.475 ;
        RECT 95.060 74.305 96.465 74.475 ;
        RECT 93.590 73.965 95.690 74.135 ;
        RECT 93.590 73.730 93.760 73.965 ;
        RECT 95.360 73.885 95.690 73.965 ;
        RECT 94.470 73.605 95.190 73.795 ;
        RECT 93.590 72.945 93.760 73.560 ;
        RECT 93.930 73.435 94.260 73.580 ;
        RECT 93.930 73.115 95.220 73.435 ;
        RECT 95.390 72.945 95.560 73.660 ;
        RECT 93.590 72.775 95.560 72.945 ;
        RECT 92.595 72.290 93.840 72.500 ;
        RECT 92.595 71.530 93.310 72.290 ;
        RECT 94.220 72.070 94.550 72.775 ;
        RECT 94.755 72.050 95.130 72.605 ;
        RECT 95.860 72.595 96.465 74.305 ;
        RECT 98.035 74.575 99.295 74.780 ;
        RECT 100.865 75.680 101.470 76.160 ;
        RECT 101.640 76.040 102.575 76.190 ;
        RECT 103.280 76.040 103.805 76.170 ;
        RECT 101.640 75.850 103.805 76.040 ;
        RECT 102.780 75.840 103.805 75.850 ;
        RECT 104.020 76.160 104.190 76.430 ;
        RECT 104.760 76.330 105.770 76.610 ;
        RECT 105.940 76.435 107.345 76.690 ;
        RECT 106.740 76.335 107.345 76.435 ;
        RECT 108.915 76.875 110.175 78.460 ;
        RECT 108.915 76.535 111.005 76.875 ;
        RECT 108.915 76.335 110.175 76.535 ;
        RECT 106.740 76.160 106.910 76.335 ;
        RECT 109.460 76.160 110.175 76.335 ;
        RECT 100.865 75.510 102.480 75.680 ;
        RECT 100.865 74.840 101.470 75.510 ;
        RECT 101.685 75.165 102.610 75.340 ;
        RECT 102.780 75.290 103.110 75.840 ;
        RECT 104.020 75.670 104.735 76.160 ;
        RECT 103.410 75.500 104.735 75.670 ;
        RECT 103.280 75.175 103.800 75.330 ;
        RECT 101.685 75.120 102.660 75.165 ;
        RECT 103.240 75.120 103.800 75.175 ;
        RECT 101.685 75.010 103.800 75.120 ;
        RECT 102.530 75.000 103.800 75.010 ;
        RECT 102.530 74.950 103.365 75.000 ;
        RECT 100.865 74.670 102.385 74.840 ;
        RECT 104.020 74.830 104.735 75.500 ;
        RECT 98.035 74.235 100.125 74.575 ;
        RECT 100.865 74.320 101.470 74.670 ;
        RECT 103.505 74.660 104.735 74.830 ;
        RECT 104.020 74.575 104.735 74.660 ;
        RECT 98.035 73.195 99.295 74.235 ;
        RECT 97.205 72.855 99.295 73.195 ;
        RECT 95.360 72.280 96.465 72.595 ;
        RECT 93.525 71.900 94.050 72.030 ;
        RECT 94.755 71.900 95.690 72.050 ;
        RECT 93.525 71.710 95.690 71.900 ;
        RECT 93.525 71.700 94.550 71.710 ;
        RECT 92.595 71.360 93.920 71.530 ;
        RECT 92.595 71.275 93.310 71.360 ;
        RECT 88.085 70.980 88.610 71.110 ;
        RECT 89.315 70.980 90.250 71.130 ;
        RECT 88.085 70.790 90.250 70.980 ;
        RECT 90.420 71.100 90.590 71.275 ;
        RECT 93.140 71.100 93.310 71.275 ;
        RECT 88.085 70.780 89.110 70.790 ;
        RECT 86.410 70.440 88.480 70.610 ;
        RECT 86.410 70.370 87.870 70.440 ;
        RECT 84.980 70.180 86.760 70.200 ;
        RECT 80.970 68.990 83.720 70.180 ;
        RECT 81.490 68.970 83.720 68.990 ;
        RECT 73.665 67.595 74.270 68.055 ;
        RECT 71.380 66.960 71.550 67.595 ;
        RECT 74.100 66.960 74.270 67.595 ;
        RECT 76.820 67.130 77.760 68.055 ;
        RECT 77.930 67.130 81.320 68.820 ;
        RECT 81.490 67.590 83.200 68.970 ;
        RECT 83.890 68.800 86.760 70.180 ;
        RECT 83.370 68.510 86.760 68.800 ;
        RECT 86.930 69.770 87.870 70.370 ;
        RECT 88.090 70.115 88.610 70.270 ;
        RECT 88.780 70.230 89.110 70.780 ;
        RECT 90.420 70.620 91.680 71.100 ;
        RECT 89.410 70.450 91.680 70.620 ;
        RECT 88.090 70.060 88.650 70.115 ;
        RECT 89.280 70.105 90.205 70.280 ;
        RECT 89.230 70.060 90.205 70.105 ;
        RECT 88.090 69.950 90.205 70.060 ;
        RECT 88.090 69.940 89.360 69.950 ;
        RECT 88.525 69.890 89.360 69.940 ;
        RECT 90.420 69.780 91.680 70.450 ;
        RECT 86.930 69.600 88.385 69.770 ;
        RECT 89.505 69.610 91.680 69.780 ;
        RECT 86.930 69.260 87.870 69.600 ;
        RECT 90.420 69.280 91.680 69.610 ;
        RECT 91.850 70.690 93.310 71.100 ;
        RECT 93.530 71.035 94.050 71.190 ;
        RECT 94.220 71.150 94.550 71.700 ;
        RECT 95.860 71.540 96.465 72.280 ;
        RECT 94.850 71.375 96.465 71.540 ;
        RECT 94.850 71.370 97.715 71.375 ;
        RECT 93.530 70.980 94.090 71.035 ;
        RECT 94.720 71.025 95.645 71.200 ;
        RECT 94.670 70.980 95.645 71.025 ;
        RECT 93.530 70.870 95.645 70.980 ;
        RECT 95.860 71.025 97.715 71.370 ;
        RECT 93.530 70.860 94.800 70.870 ;
        RECT 93.965 70.810 94.800 70.860 ;
        RECT 95.860 70.700 96.465 71.025 ;
        RECT 91.850 70.520 93.825 70.690 ;
        RECT 94.945 70.530 96.465 70.700 ;
        RECT 91.850 70.180 93.310 70.520 ;
        RECT 95.860 70.180 96.465 70.530 ;
        RECT 91.850 69.450 94.600 70.180 ;
        RECT 90.420 69.260 92.200 69.280 ;
        RECT 86.930 68.510 89.160 69.260 ;
        RECT 83.370 68.340 85.150 68.510 ;
        RECT 87.700 68.340 88.640 68.510 ;
        RECT 89.330 68.340 92.200 69.260 ;
        RECT 83.370 67.650 86.240 68.340 ;
        RECT 86.410 67.820 88.640 68.340 ;
        RECT 83.370 67.590 86.780 67.650 ;
        RECT 81.490 67.130 82.430 67.590 ;
        RECT 76.820 66.960 76.990 67.130 ;
        RECT 79.540 66.960 79.710 67.130 ;
        RECT 82.260 66.960 82.430 67.130 ;
        RECT 84.980 67.130 86.780 67.590 ;
        RECT 86.950 67.590 88.640 67.820 ;
        RECT 88.810 67.590 92.200 68.340 ;
        RECT 92.370 68.970 94.600 69.450 ;
        RECT 94.770 69.435 96.465 70.180 ;
        RECT 98.035 70.815 99.295 72.855 ;
        RECT 100.865 74.060 102.610 74.320 ;
        RECT 100.865 73.390 101.470 74.060 ;
        RECT 101.640 73.560 102.610 73.890 ;
        RECT 102.780 73.560 103.030 74.320 ;
        RECT 103.220 73.980 103.850 74.320 ;
        RECT 104.020 74.235 105.565 74.575 ;
        RECT 100.865 73.220 102.270 73.390 ;
        RECT 100.865 72.755 101.470 73.220 ;
        RECT 102.440 73.050 102.610 73.560 ;
        RECT 103.220 73.470 103.390 73.980 ;
        RECT 104.020 73.810 104.735 74.235 ;
        RECT 103.560 73.640 104.735 73.810 ;
        RECT 99.615 72.550 101.470 72.755 ;
        RECT 101.640 72.720 102.610 73.050 ;
        RECT 99.615 72.405 102.270 72.550 ;
        RECT 100.865 72.295 102.270 72.405 ;
        RECT 102.440 72.470 102.610 72.720 ;
        RECT 102.780 72.640 103.030 73.390 ;
        RECT 103.220 73.220 103.850 73.470 ;
        RECT 103.200 72.470 103.450 73.050 ;
        RECT 103.640 72.630 103.850 73.220 ;
        RECT 100.865 72.020 101.470 72.295 ;
        RECT 102.440 72.190 103.450 72.470 ;
        RECT 103.620 72.300 103.850 72.630 ;
        RECT 104.020 72.020 104.735 73.640 ;
        RECT 106.305 72.755 107.345 76.160 ;
        RECT 108.915 74.575 110.175 76.160 ;
        RECT 111.745 75.055 112.350 78.460 ;
        RECT 110.495 74.705 112.350 75.055 ;
        RECT 108.085 74.235 110.175 74.575 ;
        RECT 108.915 73.115 110.175 74.235 ;
        RECT 111.745 73.115 112.350 74.705 ;
        RECT 108.915 72.940 109.630 73.115 ;
        RECT 112.180 72.940 112.350 73.115 ;
        RECT 105.055 72.405 108.595 72.755 ;
        RECT 100.865 70.815 102.560 72.020 ;
        RECT 98.035 70.640 98.750 70.815 ;
        RECT 101.300 70.640 102.560 70.815 ;
        RECT 98.035 69.435 100.040 70.640 ;
        RECT 94.770 69.260 96.030 69.435 ;
        RECT 98.580 69.260 100.040 69.435 ;
        RECT 92.370 67.590 94.080 68.970 ;
        RECT 94.770 68.800 97.120 69.260 ;
        RECT 94.250 68.340 97.120 68.800 ;
        RECT 97.290 68.990 100.040 69.260 ;
        RECT 100.210 70.200 102.560 70.640 ;
        RECT 102.730 70.815 104.735 72.020 ;
        RECT 106.305 70.815 107.345 72.405 ;
        RECT 108.915 71.355 110.175 72.940 ;
        RECT 108.915 71.015 111.005 71.355 ;
        RECT 108.915 70.815 110.175 71.015 ;
        RECT 102.730 70.640 104.190 70.815 ;
        RECT 106.740 70.640 106.910 70.815 ;
        RECT 109.460 70.640 110.175 70.815 ;
        RECT 102.730 70.370 105.480 70.640 ;
        RECT 97.290 68.510 99.520 68.990 ;
        RECT 100.210 68.820 103.080 70.200 ;
        RECT 94.250 67.590 97.640 68.340 ;
        RECT 97.810 67.590 99.520 68.510 ;
        RECT 86.950 67.130 87.870 67.590 ;
        RECT 84.980 66.960 85.150 67.130 ;
        RECT 87.700 66.960 87.870 67.130 ;
        RECT 90.420 66.960 90.590 67.590 ;
        RECT 93.140 66.960 93.310 67.590 ;
        RECT 95.860 66.960 96.030 67.590 ;
        RECT 98.580 67.130 99.520 67.590 ;
        RECT 99.690 68.510 103.080 68.820 ;
        RECT 103.250 68.990 105.480 70.370 ;
        RECT 103.250 68.510 104.960 68.990 ;
        RECT 105.650 68.820 108.000 70.640 ;
        RECT 108.170 68.990 110.175 70.640 ;
        RECT 111.745 69.535 112.350 72.940 ;
        RECT 110.495 69.185 112.350 69.535 ;
        RECT 99.690 68.340 101.470 68.510 ;
        RECT 104.020 68.340 104.960 68.510 ;
        RECT 99.690 67.650 102.560 68.340 ;
        RECT 102.730 67.820 104.960 68.340 ;
        RECT 99.690 67.130 103.100 67.650 ;
        RECT 103.270 67.130 104.960 67.820 ;
        RECT 105.130 67.130 108.520 68.820 ;
        RECT 108.690 67.595 110.175 68.990 ;
        RECT 111.745 67.595 112.350 69.185 ;
        RECT 108.690 67.130 109.630 67.595 ;
        RECT 98.580 66.960 98.750 67.130 ;
        RECT 101.300 66.960 101.470 67.130 ;
        RECT 104.020 66.960 104.190 67.130 ;
        RECT 106.740 66.960 106.910 67.130 ;
        RECT 109.460 66.960 109.630 67.130 ;
        RECT 112.180 66.960 112.350 67.595 ;
        RECT 60.500 66.270 61.420 66.960 ;
        RECT 61.590 66.440 65.020 66.960 ;
        RECT 60.500 65.750 61.960 66.270 ;
        RECT 62.130 65.750 64.480 66.440 ;
        RECT 65.190 66.270 66.860 66.960 ;
        RECT 67.030 66.440 70.460 66.960 ;
        RECT 64.650 65.750 67.400 66.270 ;
        RECT 67.570 65.750 69.920 66.440 ;
        RECT 70.630 66.270 72.300 66.960 ;
        RECT 72.470 66.440 75.900 66.960 ;
        RECT 70.090 65.750 72.840 66.270 ;
        RECT 73.010 65.750 75.360 66.440 ;
        RECT 76.070 66.270 77.740 66.960 ;
        RECT 77.910 66.440 81.340 66.960 ;
        RECT 75.530 65.750 78.280 66.270 ;
        RECT 78.450 65.750 80.800 66.440 ;
        RECT 81.510 66.270 83.180 66.960 ;
        RECT 83.350 66.440 86.780 66.960 ;
        RECT 80.970 65.750 83.720 66.270 ;
        RECT 83.890 65.750 86.240 66.440 ;
        RECT 86.950 66.270 88.620 66.960 ;
        RECT 88.790 66.440 92.220 66.960 ;
        RECT 86.410 65.750 89.160 66.270 ;
        RECT 89.330 65.750 91.680 66.440 ;
        RECT 92.390 66.270 94.060 66.960 ;
        RECT 94.230 66.440 97.660 66.960 ;
        RECT 91.850 65.750 94.600 66.270 ;
        RECT 94.770 65.750 97.120 66.440 ;
        RECT 97.830 66.270 99.500 66.960 ;
        RECT 99.670 66.440 103.100 66.960 ;
        RECT 97.290 65.750 100.040 66.270 ;
        RECT 100.210 65.750 102.560 66.440 ;
        RECT 103.270 66.270 104.940 66.960 ;
        RECT 105.110 66.440 108.540 66.960 ;
        RECT 102.730 65.750 105.480 66.270 ;
        RECT 105.650 65.750 108.000 66.440 ;
        RECT 108.710 66.270 110.380 66.960 ;
        RECT 110.550 66.440 112.350 66.960 ;
        RECT 108.170 65.750 110.920 66.270 ;
        RECT 111.090 65.750 112.350 66.440 ;
        RECT 60.500 65.665 60.670 65.750 ;
        RECT 63.220 65.665 63.390 65.750 ;
        RECT 65.940 65.665 66.110 65.750 ;
        RECT 68.660 65.665 68.830 65.750 ;
        RECT 71.380 65.665 71.550 65.750 ;
        RECT 74.100 65.665 74.270 65.750 ;
        RECT 76.820 65.665 76.990 65.750 ;
        RECT 79.540 65.665 79.710 65.750 ;
        RECT 82.260 65.665 82.430 65.750 ;
        RECT 84.980 65.665 85.150 65.750 ;
        RECT 87.700 65.665 87.870 65.750 ;
        RECT 90.420 65.665 90.590 65.750 ;
        RECT 93.140 65.665 93.310 65.750 ;
        RECT 95.860 65.665 96.030 65.750 ;
        RECT 98.580 65.665 98.750 65.750 ;
        RECT 101.300 65.665 101.470 65.750 ;
        RECT 104.020 65.665 104.190 65.750 ;
        RECT 106.740 65.665 106.910 65.750 ;
        RECT 109.460 65.665 109.630 65.750 ;
        RECT 112.180 65.665 112.350 65.750 ;
        RECT 13.525 21.570 13.875 21.970 ;
        RECT 17.120 21.575 17.495 21.970 ;
        RECT 12.425 19.180 12.825 21.570 ;
        RECT 13.075 19.770 13.875 21.570 ;
        RECT 16.045 19.265 16.445 21.575 ;
        RECT 16.695 19.775 17.495 21.575 ;
        RECT 13.275 19.180 13.600 19.230 ;
        RECT 12.425 18.980 13.600 19.180 ;
        RECT 12.425 18.260 12.825 18.980 ;
        RECT 13.275 18.905 13.600 18.980 ;
        RECT 15.970 18.670 16.565 19.265 ;
        RECT 12.425 17.800 12.905 18.260 ;
        RECT 12.505 17.460 12.905 17.800 ;
        RECT 13.155 17.460 13.955 18.260 ;
        RECT 16.045 18.255 16.445 18.670 ;
        RECT 16.045 17.710 16.530 18.255 ;
        RECT 13.555 16.985 13.955 17.460 ;
        RECT 16.130 17.455 16.530 17.710 ;
        RECT 16.780 17.455 17.580 18.255 ;
        RECT 17.180 16.985 17.580 17.455 ;
        RECT 12.605 16.205 13.200 16.800 ;
        RECT 13.555 16.725 17.580 16.985 ;
        RECT 14.250 15.990 14.845 16.585 ;
        RECT 13.870 14.920 14.670 15.720 ;
        RECT 14.920 14.920 15.320 16.725 ;
        RECT 16.325 15.680 16.930 16.180 ;
        RECT 13.870 14.370 14.270 14.920 ;
        RECT 12.885 12.645 13.685 13.995 ;
        RECT 13.935 12.595 14.335 13.445 ;
        RECT 15.135 13.430 15.940 13.995 ;
        RECT 15.140 12.640 15.940 13.430 ;
        RECT 13.960 12.525 14.335 12.595 ;
        RECT 16.190 12.575 16.590 13.440 ;
        RECT 17.390 12.650 18.190 14.000 ;
        RECT 18.440 12.595 18.840 13.450 ;
        RECT 19.645 12.645 20.445 13.995 ;
        RECT 20.695 12.600 21.095 13.445 ;
        RECT 20.705 12.595 21.095 12.600 ;
        RECT 14.035 12.425 14.335 12.525 ;
        RECT 16.330 12.425 16.590 12.575 ;
        RECT 18.460 12.525 18.840 12.595 ;
        RECT 18.485 12.430 18.840 12.525 ;
        RECT 14.035 12.405 16.020 12.425 ;
        RECT 13.420 11.955 13.825 12.250 ;
        RECT 14.035 12.125 16.085 12.405 ;
        RECT 16.330 12.195 18.290 12.425 ;
        RECT 16.330 12.130 18.270 12.195 ;
        RECT 9.710 10.965 10.110 11.515 ;
        RECT 8.660 10.165 9.060 10.965 ;
        RECT 9.310 10.165 10.110 10.965 ;
        RECT 13.435 10.275 13.835 10.675 ;
        RECT 8.660 9.865 8.910 10.165 ;
        RECT 14.035 10.075 14.335 12.125 ;
        RECT 15.735 10.775 16.135 11.130 ;
        RECT 16.330 10.575 16.590 12.130 ;
        RECT 17.885 12.025 18.270 12.130 ;
        RECT 18.485 12.145 20.535 12.430 ;
        RECT 18.485 12.120 20.525 12.145 ;
        RECT 18.485 12.025 18.840 12.120 ;
        RECT 9.110 9.765 10.310 9.865 ;
        RECT 9.110 9.565 10.060 9.765 ;
        RECT 10.260 9.565 10.310 9.765 ;
        RECT 9.110 9.465 10.310 9.565 ;
        RECT 8.660 8.965 8.910 9.465 ;
        RECT 8.660 8.165 9.060 8.965 ;
        RECT 9.310 8.165 10.110 8.965 ;
        RECT 8.660 7.165 9.060 7.965 ;
        RECT 9.310 7.165 10.110 7.965 ;
        RECT 9.710 6.765 10.110 7.165 ;
        RECT 12.885 6.770 13.685 8.965 ;
        RECT 13.935 7.165 14.335 10.075 ;
        RECT 15.140 6.760 15.940 8.960 ;
        RECT 16.190 7.160 16.590 10.575 ;
        RECT 18.440 9.800 18.840 12.025 ;
        RECT 20.735 11.975 21.095 12.595 ;
        RECT 20.695 10.325 21.095 11.975 ;
        RECT 77.675 12.950 78.075 13.350 ;
        RECT 18.455 9.725 18.840 9.800 ;
        RECT 20.085 9.780 20.585 10.120 ;
        RECT 20.785 9.865 21.095 10.325 ;
        RECT 23.655 10.965 24.055 11.515 ;
        RECT 77.675 11.150 78.475 12.950 ;
        RECT 78.725 11.150 79.125 12.950 ;
        RECT 23.655 10.165 24.455 10.965 ;
        RECT 24.705 10.165 25.105 10.965 ;
        RECT 78.875 10.650 79.125 11.150 ;
        RECT 80.825 11.055 81.625 12.950 ;
        RECT 81.875 11.150 82.275 12.950 ;
        RECT 80.825 10.805 81.225 11.055 ;
        RECT 77.525 10.350 77.725 10.550 ;
        RECT 78.275 10.250 78.675 10.650 ;
        RECT 78.875 10.250 79.325 10.650 ;
        RECT 79.605 10.585 81.225 10.805 ;
        RECT 24.855 9.865 25.105 10.165 ;
        RECT 78.875 9.950 79.125 10.250 ;
        RECT 17.775 9.295 18.285 9.630 ;
        RECT 17.775 9.220 18.270 9.295 ;
        RECT 18.485 9.125 18.840 9.725 ;
        RECT 20.785 9.765 24.655 9.865 ;
        RECT 20.785 9.570 23.505 9.765 ;
        RECT 17.380 6.770 18.190 8.970 ;
        RECT 18.440 7.170 18.840 9.125 ;
        RECT 20.695 9.565 23.505 9.570 ;
        RECT 23.705 9.565 24.655 9.765 ;
        RECT 20.695 9.465 24.655 9.565 ;
        RECT 19.645 6.765 20.445 8.965 ;
        RECT 20.695 7.165 21.095 9.465 ;
        RECT 24.855 8.965 25.105 9.465 ;
        RECT 23.655 8.165 24.455 8.965 ;
        RECT 24.705 8.165 25.105 8.965 ;
        RECT 77.675 9.150 78.475 9.950 ;
        RECT 78.725 9.150 79.125 9.950 ;
        RECT 77.675 8.600 78.075 9.150 ;
        RECT 79.605 9.050 79.855 10.585 ;
        RECT 80.025 9.650 80.425 10.055 ;
        RECT 80.825 9.950 81.225 10.585 ;
        RECT 81.630 10.555 81.800 10.725 ;
        RECT 82.025 10.650 82.275 11.150 ;
        RECT 82.025 10.250 82.475 10.650 ;
        RECT 82.025 9.950 82.275 10.250 ;
        RECT 80.825 9.150 81.625 9.950 ;
        RECT 81.875 9.150 82.275 9.950 ;
        RECT 79.605 8.610 80.165 9.050 ;
        RECT 23.655 7.165 24.455 7.965 ;
        RECT 24.705 7.165 25.105 7.965 ;
        RECT 23.655 6.765 24.055 7.165 ;
      LAYER met1 ;
        RECT 55.485 213.020 55.785 225.755 ;
        RECT 16.590 213.015 55.785 213.020 ;
        RECT 16.565 212.520 55.785 213.015 ;
        RECT 16.565 204.495 16.960 212.520 ;
        RECT 58.260 212.025 58.590 225.765 ;
        RECT 61.030 225.465 61.290 225.765 ;
        RECT 63.800 225.480 64.080 225.760 ;
        RECT 61.015 225.185 61.295 225.465 ;
        RECT 63.785 225.200 64.080 225.480 ;
        RECT 19.685 212.015 58.590 212.025 ;
        RECT 19.680 211.720 58.590 212.015 ;
        RECT 19.680 204.640 20.035 211.720 ;
        RECT 61.030 210.995 61.290 225.185 ;
        RECT 23.380 210.740 61.290 210.995 ;
        RECT 16.565 204.145 16.965 204.495 ;
        RECT 19.665 204.345 20.175 204.640 ;
        RECT 23.380 204.580 23.695 210.740 ;
        RECT 28.170 210.120 28.480 210.125 ;
        RECT 63.800 210.120 64.080 225.200 ;
        RECT 28.170 209.920 64.080 210.120 ;
        RECT 28.170 209.915 63.625 209.920 ;
        RECT 28.170 204.700 28.480 209.915 ;
        RECT 32.355 208.975 32.740 209.005 ;
        RECT 66.505 208.975 66.920 225.775 ;
        RECT 32.355 208.530 66.920 208.975 ;
        RECT 69.300 225.515 69.605 225.765 ;
        RECT 69.300 225.235 69.610 225.515 ;
        RECT 23.365 204.195 24.120 204.580 ;
        RECT 28.165 204.395 28.760 204.700 ;
        RECT 32.355 204.595 32.740 208.530 ;
        RECT 53.020 207.750 53.455 207.760 ;
        RECT 69.300 207.750 69.605 225.235 ;
        RECT 53.020 207.415 69.605 207.750 ;
        RECT 32.355 204.480 33.115 204.595 ;
        RECT 32.365 204.195 33.115 204.480 ;
        RECT 48.995 203.820 50.500 204.000 ;
        RECT 16.410 203.520 50.500 203.820 ;
        RECT 18.210 203.515 50.500 203.520 ;
        RECT 48.995 203.310 50.500 203.515 ;
        RECT 1.000 198.855 2.500 199.255 ;
        RECT 1.000 198.560 17.860 198.855 ;
        RECT 1.000 198.240 2.500 198.560 ;
        RECT 15.625 198.555 17.860 198.560 ;
        RECT 19.065 198.850 20.700 198.855 ;
        RECT 19.065 198.570 21.470 198.850 ;
        RECT 19.065 198.555 21.475 198.570 ;
        RECT 21.120 196.770 21.475 198.555 ;
        RECT 21.120 196.470 25.865 196.770 ;
        RECT 25.500 192.900 25.865 196.470 ;
        RECT 25.500 192.600 30.565 192.900 ;
        RECT 30.360 185.030 30.565 192.600 ;
        RECT 30.360 184.905 33.210 185.030 ;
        RECT 30.360 184.730 33.465 184.905 ;
        RECT 30.820 38.960 31.135 184.730 ;
        RECT 53.020 46.155 53.455 207.415 ;
        RECT 60.345 65.665 60.825 117.645 ;
        RECT 61.645 114.035 61.905 114.355 ;
        RECT 61.705 112.140 61.845 114.035 ;
        RECT 61.985 113.115 62.245 113.435 ;
        RECT 62.340 112.645 62.570 112.935 ;
        RECT 62.000 112.250 62.230 112.540 ;
        RECT 61.660 111.850 61.890 112.140 ;
        RECT 62.045 111.350 62.185 112.250 ;
        RECT 62.000 111.060 62.230 111.350 ;
        RECT 62.045 108.830 62.185 111.060 ;
        RECT 62.385 110.835 62.525 112.645 ;
        RECT 62.340 110.545 62.570 110.835 ;
        RECT 62.385 109.265 62.525 110.545 ;
        RECT 62.340 108.975 62.570 109.265 ;
        RECT 62.000 108.540 62.230 108.830 ;
        RECT 62.665 106.215 62.925 106.535 ;
        RECT 62.725 102.855 62.865 106.215 ;
        RECT 62.665 102.535 62.925 102.855 ;
        RECT 61.645 99.775 61.905 100.095 ;
        RECT 61.705 97.780 61.845 99.775 ;
        RECT 61.660 97.490 61.890 97.780 ;
        RECT 61.645 97.015 61.905 97.335 ;
        RECT 62.680 97.030 62.910 97.320 ;
        RECT 61.705 96.860 61.845 97.015 ;
        RECT 61.660 96.570 61.890 96.860 ;
        RECT 61.705 90.880 61.845 96.570 ;
        RECT 62.725 96.415 62.865 97.030 ;
        RECT 62.665 96.095 62.925 96.415 ;
        RECT 61.985 93.335 62.245 93.655 ;
        RECT 62.045 91.340 62.185 93.335 ;
        RECT 62.000 91.050 62.230 91.340 ;
        RECT 61.660 90.805 61.890 90.880 ;
        RECT 61.660 90.665 62.185 90.805 ;
        RECT 61.660 90.590 61.890 90.665 ;
        RECT 61.645 90.115 61.905 90.435 ;
        RECT 61.705 89.960 61.845 90.115 ;
        RECT 61.660 89.670 61.890 89.960 ;
        RECT 62.045 82.155 62.185 90.665 ;
        RECT 61.985 81.835 62.245 82.155 ;
        RECT 62.340 80.470 62.570 80.760 ;
        RECT 62.385 75.255 62.525 80.470 ;
        RECT 62.665 79.995 62.925 80.315 ;
        RECT 62.725 79.840 62.865 79.995 ;
        RECT 62.680 79.550 62.910 79.840 ;
        RECT 62.325 74.935 62.585 75.255 ;
        RECT 63.065 65.665 63.545 117.645 ;
        RECT 64.705 113.345 64.965 113.435 ;
        RECT 64.705 113.205 65.585 113.345 ;
        RECT 64.705 113.115 64.965 113.205 ;
        RECT 64.040 112.645 64.270 112.935 ;
        RECT 65.045 112.655 65.305 112.975 ;
        RECT 64.085 110.835 64.225 112.645 ;
        RECT 64.380 112.250 64.610 112.540 ;
        RECT 64.425 111.350 64.565 112.250 ;
        RECT 65.105 112.085 65.245 112.655 ;
        RECT 65.445 112.515 65.585 113.205 ;
        RECT 65.385 112.195 65.645 112.515 ;
        RECT 65.060 111.795 65.290 112.085 ;
        RECT 64.380 111.060 64.610 111.350 ;
        RECT 64.040 110.545 64.270 110.835 ;
        RECT 64.085 109.265 64.225 110.545 ;
        RECT 64.040 108.975 64.270 109.265 ;
        RECT 64.425 108.830 64.565 111.060 ;
        RECT 64.380 108.540 64.610 108.830 ;
        RECT 64.040 106.230 64.270 106.520 ;
        RECT 64.085 103.775 64.225 106.230 ;
        RECT 64.025 103.455 64.285 103.775 ;
        RECT 65.060 103.470 65.290 103.760 ;
        RECT 64.720 102.765 64.950 102.840 ;
        RECT 63.745 102.625 64.950 102.765 ;
        RECT 63.745 97.335 63.885 102.625 ;
        RECT 64.720 102.550 64.950 102.625 ;
        RECT 65.105 102.395 65.245 103.470 ;
        RECT 64.365 102.075 64.625 102.395 ;
        RECT 65.045 102.075 65.305 102.395 ;
        RECT 63.685 97.245 63.945 97.335 ;
        RECT 64.425 97.320 64.565 102.075 ;
        RECT 65.060 101.630 65.290 101.920 ;
        RECT 65.105 100.095 65.245 101.630 ;
        RECT 65.045 99.775 65.305 100.095 ;
        RECT 64.720 99.330 64.950 99.620 ;
        RECT 63.685 97.105 64.225 97.245 ;
        RECT 63.685 97.015 63.945 97.105 ;
        RECT 63.700 96.570 63.930 96.860 ;
        RECT 63.745 95.940 63.885 96.570 ;
        RECT 63.700 95.650 63.930 95.940 ;
        RECT 64.085 94.945 64.225 97.105 ;
        RECT 64.380 97.030 64.610 97.320 ;
        RECT 64.425 95.955 64.565 97.030 ;
        RECT 64.765 96.860 64.905 99.330 ;
        RECT 64.720 96.785 64.950 96.860 ;
        RECT 64.720 96.645 65.245 96.785 ;
        RECT 64.720 96.570 64.950 96.645 ;
        RECT 64.365 95.635 64.625 95.955 ;
        RECT 64.085 94.805 64.905 94.945 ;
        RECT 64.365 94.255 64.625 94.575 ;
        RECT 64.025 93.795 64.285 94.115 ;
        RECT 64.040 88.725 64.270 89.015 ;
        RECT 64.425 88.965 64.565 94.255 ;
        RECT 64.765 93.180 64.905 94.805 ;
        RECT 64.720 92.890 64.950 93.180 ;
        RECT 65.105 92.260 65.245 96.645 ;
        RECT 65.060 91.970 65.290 92.260 ;
        RECT 65.105 90.895 65.245 91.970 ;
        RECT 65.045 90.575 65.305 90.895 ;
        RECT 64.720 89.425 64.950 89.500 ;
        RECT 65.445 89.425 65.585 112.195 ;
        RECT 64.720 89.285 65.585 89.425 ;
        RECT 64.720 89.210 64.950 89.285 ;
        RECT 64.425 88.825 64.905 88.965 ;
        RECT 64.085 86.915 64.225 88.725 ;
        RECT 64.380 88.330 64.610 88.620 ;
        RECT 64.425 87.430 64.565 88.330 ;
        RECT 64.765 88.220 64.905 88.825 ;
        RECT 64.720 87.930 64.950 88.220 ;
        RECT 65.105 88.045 65.245 89.285 ;
        RECT 65.385 88.045 65.645 88.135 ;
        RECT 65.105 87.905 65.645 88.045 ;
        RECT 64.380 87.140 64.610 87.430 ;
        RECT 64.040 86.625 64.270 86.915 ;
        RECT 64.085 85.345 64.225 86.625 ;
        RECT 64.040 85.055 64.270 85.345 ;
        RECT 64.425 84.910 64.565 87.140 ;
        RECT 64.380 84.620 64.610 84.910 ;
        RECT 63.685 81.835 63.945 82.155 ;
        RECT 63.745 74.780 63.885 81.835 ;
        RECT 64.720 81.605 64.950 81.680 ;
        RECT 65.105 81.605 65.245 87.905 ;
        RECT 65.385 87.815 65.645 87.905 ;
        RECT 65.385 82.755 65.645 83.075 ;
        RECT 65.445 82.600 65.585 82.755 ;
        RECT 65.400 82.310 65.630 82.600 ;
        RECT 64.720 81.465 65.245 81.605 ;
        RECT 64.720 81.390 64.950 81.465 ;
        RECT 64.040 80.905 64.270 81.195 ;
        RECT 64.085 79.095 64.225 80.905 ;
        RECT 64.380 80.510 64.610 80.800 ;
        RECT 64.425 79.610 64.565 80.510 ;
        RECT 64.720 80.315 64.950 80.345 ;
        RECT 64.705 79.995 64.965 80.315 ;
        RECT 64.380 79.320 64.610 79.610 ;
        RECT 64.040 78.805 64.270 79.095 ;
        RECT 64.085 77.525 64.225 78.805 ;
        RECT 64.040 77.235 64.270 77.525 ;
        RECT 64.425 77.090 64.565 79.320 ;
        RECT 64.380 76.800 64.610 77.090 ;
        RECT 63.700 74.490 63.930 74.780 ;
        RECT 65.785 65.665 66.265 117.645 ;
        RECT 67.085 113.575 67.345 113.895 ;
        RECT 66.405 112.655 66.665 112.975 ;
        RECT 67.085 112.195 67.345 112.515 ;
        RECT 67.780 111.725 68.010 112.015 ;
        RECT 67.440 111.330 67.670 111.620 ;
        RECT 67.145 111.165 67.285 111.330 ;
        RECT 67.100 111.135 67.330 111.165 ;
        RECT 67.085 110.815 67.345 111.135 ;
        RECT 67.485 110.430 67.625 111.330 ;
        RECT 67.440 110.140 67.670 110.430 ;
        RECT 67.485 107.910 67.625 110.140 ;
        RECT 67.825 109.915 67.965 111.725 ;
        RECT 67.780 109.625 68.010 109.915 ;
        RECT 67.825 108.345 67.965 109.625 ;
        RECT 67.780 108.055 68.010 108.345 ;
        RECT 67.440 107.620 67.670 107.910 ;
        RECT 68.105 106.215 68.365 106.535 ;
        RECT 67.780 105.310 68.010 105.600 ;
        RECT 67.425 103.455 67.685 103.775 ;
        RECT 66.760 103.010 66.990 103.300 ;
        RECT 66.805 102.855 66.945 103.010 ;
        RECT 66.745 102.535 67.005 102.855 ;
        RECT 67.485 102.840 67.625 103.455 ;
        RECT 67.440 102.550 67.670 102.840 ;
        RECT 66.745 102.075 67.005 102.395 ;
        RECT 66.805 98.240 66.945 102.075 ;
        RECT 67.100 101.845 67.330 101.920 ;
        RECT 67.825 101.845 67.965 105.310 ;
        RECT 68.165 103.300 68.305 106.215 ;
        RECT 68.120 103.010 68.350 103.300 ;
        RECT 67.100 101.705 67.965 101.845 ;
        RECT 67.100 101.630 67.330 101.705 ;
        RECT 67.145 98.625 67.285 101.630 ;
        RECT 68.120 100.710 68.350 101.000 ;
        RECT 68.165 100.095 68.305 100.710 ;
        RECT 68.105 99.775 68.365 100.095 ;
        RECT 67.425 98.625 67.685 98.715 ;
        RECT 67.145 98.485 67.685 98.625 ;
        RECT 67.425 98.395 67.685 98.485 ;
        RECT 66.760 97.950 66.990 98.240 ;
        RECT 66.420 97.490 66.650 97.780 ;
        RECT 66.465 96.415 66.605 97.490 ;
        RECT 66.405 96.095 66.665 96.415 ;
        RECT 68.120 95.650 68.350 95.940 ;
        RECT 67.425 95.175 67.685 95.495 ;
        RECT 66.405 94.255 66.665 94.575 ;
        RECT 66.405 93.795 66.665 94.115 ;
        RECT 66.465 93.640 66.605 93.795 ;
        RECT 66.420 93.350 66.650 93.640 ;
        RECT 66.745 92.415 67.005 92.735 ;
        RECT 67.100 91.265 67.330 91.340 ;
        RECT 67.485 91.265 67.625 95.175 ;
        RECT 68.165 94.575 68.305 95.650 ;
        RECT 68.105 94.255 68.365 94.575 ;
        RECT 68.105 93.335 68.365 93.655 ;
        RECT 67.100 91.125 67.625 91.265 ;
        RECT 67.100 91.050 67.330 91.125 ;
        RECT 67.085 90.805 67.345 90.895 ;
        RECT 66.805 90.665 67.345 90.805 ;
        RECT 66.805 88.580 66.945 90.665 ;
        RECT 67.085 90.575 67.345 90.665 ;
        RECT 67.100 88.750 67.330 89.040 ;
        RECT 66.760 88.290 66.990 88.580 ;
        RECT 66.420 87.830 66.650 88.120 ;
        RECT 66.465 87.675 66.605 87.830 ;
        RECT 66.405 87.355 66.665 87.675 ;
        RECT 66.465 83.905 66.605 87.355 ;
        RECT 66.805 84.825 66.945 88.290 ;
        RECT 67.145 87.675 67.285 88.750 ;
        RECT 67.485 88.735 67.625 91.125 ;
        RECT 68.120 89.210 68.350 89.500 ;
        RECT 67.765 88.735 68.025 89.055 ;
        RECT 67.485 88.595 67.965 88.735 ;
        RECT 67.085 87.355 67.345 87.675 ;
        RECT 67.100 87.125 67.330 87.200 ;
        RECT 67.485 87.125 67.625 88.595 ;
        RECT 68.165 87.215 68.305 89.210 ;
        RECT 67.100 86.985 67.625 87.125 ;
        RECT 67.100 86.910 67.330 86.985 ;
        RECT 66.805 84.685 67.285 84.825 ;
        RECT 66.760 83.905 66.990 83.980 ;
        RECT 66.465 83.765 66.990 83.905 ;
        RECT 66.465 82.615 66.605 83.765 ;
        RECT 66.760 83.690 66.990 83.765 ;
        RECT 66.745 83.215 67.005 83.535 ;
        RECT 66.405 82.295 66.665 82.615 ;
        RECT 66.805 82.140 66.945 83.215 ;
        RECT 67.145 83.075 67.285 84.685 ;
        RECT 67.085 82.755 67.345 83.075 ;
        RECT 67.100 82.525 67.330 82.600 ;
        RECT 67.485 82.525 67.625 86.985 ;
        RECT 68.105 86.895 68.365 87.215 ;
        RECT 68.120 85.990 68.350 86.280 ;
        RECT 68.165 85.375 68.305 85.990 ;
        RECT 68.105 85.055 68.365 85.375 ;
        RECT 67.100 82.385 67.625 82.525 ;
        RECT 67.100 82.310 67.330 82.385 ;
        RECT 66.760 81.850 66.990 82.140 ;
        RECT 67.145 81.695 67.285 82.310 ;
        RECT 67.085 81.375 67.345 81.695 ;
        RECT 68.120 80.930 68.350 81.220 ;
        RECT 68.165 80.315 68.305 80.930 ;
        RECT 68.105 79.995 68.365 80.315 ;
        RECT 68.505 65.665 68.985 117.645 ;
        RECT 69.805 114.955 70.065 115.275 ;
        RECT 69.125 114.725 69.385 114.815 ;
        RECT 69.125 114.585 69.665 114.725 ;
        RECT 69.125 114.495 69.385 114.585 ;
        RECT 69.525 111.505 69.665 114.585 ;
        RECT 69.865 114.340 70.005 114.955 ;
        RECT 70.160 114.510 70.390 114.800 ;
        RECT 69.820 114.050 70.050 114.340 ;
        RECT 70.205 113.895 70.345 114.510 ;
        RECT 70.145 113.575 70.405 113.895 ;
        RECT 70.145 113.115 70.405 113.435 ;
        RECT 70.840 112.210 71.070 112.500 ;
        RECT 70.885 112.055 71.025 112.210 ;
        RECT 70.825 111.735 71.085 112.055 ;
        RECT 70.160 111.505 70.390 111.580 ;
        RECT 69.525 111.365 70.390 111.505 ;
        RECT 70.160 111.290 70.390 111.365 ;
        RECT 69.125 110.815 69.385 111.135 ;
        RECT 69.185 110.660 69.325 110.815 ;
        RECT 69.140 110.370 69.370 110.660 ;
        RECT 70.145 106.215 70.405 106.535 ;
        RECT 70.205 105.600 70.345 106.215 ;
        RECT 70.160 105.310 70.390 105.600 ;
        RECT 69.820 104.605 70.050 104.680 ;
        RECT 69.525 104.465 70.050 104.605 ;
        RECT 69.140 103.930 69.370 104.220 ;
        RECT 69.185 99.175 69.325 103.930 ;
        RECT 69.125 98.855 69.385 99.175 ;
        RECT 69.525 98.715 69.665 104.465 ;
        RECT 69.820 104.390 70.050 104.465 ;
        RECT 70.145 103.455 70.405 103.775 ;
        RECT 69.820 103.010 70.050 103.300 ;
        RECT 70.205 103.225 70.345 103.455 ;
        RECT 70.205 103.085 70.685 103.225 ;
        RECT 69.865 99.545 70.005 103.010 ;
        RECT 70.145 102.535 70.405 102.855 ;
        RECT 70.160 100.715 70.390 101.005 ;
        RECT 70.205 100.555 70.345 100.715 ;
        RECT 70.145 100.235 70.405 100.555 ;
        RECT 70.145 99.775 70.405 100.095 ;
        RECT 69.865 99.405 70.345 99.545 ;
        RECT 69.465 98.395 69.725 98.715 ;
        RECT 69.125 95.635 69.385 95.955 ;
        RECT 69.185 95.020 69.325 95.635 ;
        RECT 69.140 94.730 69.370 95.020 ;
        RECT 69.525 94.485 69.665 98.395 ;
        RECT 69.805 97.935 70.065 98.255 ;
        RECT 70.205 97.320 70.345 99.405 ;
        RECT 70.160 97.030 70.390 97.320 ;
        RECT 70.205 95.955 70.345 97.030 ;
        RECT 70.145 95.635 70.405 95.955 ;
        RECT 69.805 95.175 70.065 95.495 ;
        RECT 70.545 95.405 70.685 103.085 ;
        RECT 70.825 96.095 71.085 96.415 ;
        RECT 70.885 95.940 71.025 96.095 ;
        RECT 70.840 95.650 71.070 95.940 ;
        RECT 70.205 95.265 70.685 95.405 ;
        RECT 70.205 95.020 70.345 95.265 ;
        RECT 70.825 95.175 71.085 95.495 ;
        RECT 70.160 94.730 70.390 95.020 ;
        RECT 69.820 94.485 70.050 94.560 ;
        RECT 69.525 94.345 70.050 94.485 ;
        RECT 69.820 94.270 70.050 94.345 ;
        RECT 70.885 93.180 71.025 95.175 ;
        RECT 70.840 92.890 71.070 93.180 ;
        RECT 70.885 89.975 71.025 92.890 ;
        RECT 70.160 89.885 70.390 89.960 ;
        RECT 70.160 89.745 70.685 89.885 ;
        RECT 70.160 89.670 70.390 89.745 ;
        RECT 69.480 89.185 69.710 89.475 ;
        RECT 69.525 87.375 69.665 89.185 ;
        RECT 69.820 88.790 70.050 89.080 ;
        RECT 69.865 87.890 70.005 88.790 ;
        RECT 70.160 88.335 70.390 88.625 ;
        RECT 69.820 87.600 70.050 87.890 ;
        RECT 69.480 87.085 69.710 87.375 ;
        RECT 69.525 85.805 69.665 87.085 ;
        RECT 69.480 85.515 69.710 85.805 ;
        RECT 69.865 85.370 70.005 87.600 ;
        RECT 70.205 86.295 70.345 88.335 ;
        RECT 70.545 88.135 70.685 89.745 ;
        RECT 70.825 89.655 71.085 89.975 ;
        RECT 70.485 87.815 70.745 88.135 ;
        RECT 70.145 85.975 70.405 86.295 ;
        RECT 69.820 85.080 70.050 85.370 ;
        RECT 69.465 83.215 69.725 83.535 ;
        RECT 69.525 81.680 69.665 83.215 ;
        RECT 70.145 82.065 70.405 82.155 ;
        RECT 70.545 82.065 70.685 87.815 ;
        RECT 70.840 82.770 71.070 83.060 ;
        RECT 70.145 81.925 70.685 82.065 ;
        RECT 70.145 81.835 70.405 81.925 ;
        RECT 69.480 81.390 69.710 81.680 ;
        RECT 69.820 79.080 70.050 79.370 ;
        RECT 69.480 78.645 69.710 78.935 ;
        RECT 69.525 77.365 69.665 78.645 ;
        RECT 69.480 77.075 69.710 77.365 ;
        RECT 69.125 75.855 69.385 76.175 ;
        RECT 69.185 74.705 69.325 75.855 ;
        RECT 69.525 75.265 69.665 77.075 ;
        RECT 69.865 76.850 70.005 79.080 ;
        RECT 70.205 77.005 70.345 81.835 ;
        RECT 70.885 81.695 71.025 82.770 ;
        RECT 70.825 81.375 71.085 81.695 ;
        RECT 70.825 80.915 71.085 81.235 ;
        RECT 70.205 76.865 70.685 77.005 ;
        RECT 69.820 76.560 70.050 76.850 ;
        RECT 69.865 75.660 70.005 76.560 ;
        RECT 70.205 76.175 70.345 76.325 ;
        RECT 70.145 75.855 70.405 76.175 ;
        RECT 70.160 75.825 70.390 75.855 ;
        RECT 69.820 75.370 70.050 75.660 ;
        RECT 70.545 75.625 70.685 76.865 ;
        RECT 70.205 75.485 70.685 75.625 ;
        RECT 69.480 74.975 69.710 75.265 ;
        RECT 70.205 74.780 70.345 75.485 ;
        RECT 70.485 74.935 70.745 75.255 ;
        RECT 69.185 74.565 69.665 74.705 ;
        RECT 69.125 73.095 69.385 73.415 ;
        RECT 69.525 72.480 69.665 74.565 ;
        RECT 70.160 74.490 70.390 74.780 ;
        RECT 70.545 74.320 70.685 74.935 ;
        RECT 70.500 74.030 70.730 74.320 ;
        RECT 70.885 73.400 71.025 80.915 ;
        RECT 70.840 73.110 71.070 73.400 ;
        RECT 69.480 72.190 69.710 72.480 ;
        RECT 71.225 65.665 71.705 117.645 ;
        RECT 72.525 114.955 72.785 115.275 ;
        RECT 72.200 114.050 72.430 114.340 ;
        RECT 72.245 111.275 72.385 114.050 ;
        RECT 72.525 112.655 72.785 112.975 ;
        RECT 72.525 112.195 72.785 112.515 ;
        RECT 73.220 111.725 73.450 112.015 ;
        RECT 72.880 111.330 73.110 111.620 ;
        RECT 72.200 110.985 72.430 111.275 ;
        RECT 72.925 110.430 73.065 111.330 ;
        RECT 72.880 110.140 73.110 110.430 ;
        RECT 72.925 107.910 73.065 110.140 ;
        RECT 73.265 109.915 73.405 111.725 ;
        RECT 73.220 109.625 73.450 109.915 ;
        RECT 73.265 108.345 73.405 109.625 ;
        RECT 73.220 108.055 73.450 108.345 ;
        RECT 72.880 107.620 73.110 107.910 ;
        RECT 71.860 105.310 72.090 105.600 ;
        RECT 71.905 102.855 72.045 105.310 ;
        RECT 71.845 102.535 72.105 102.855 ;
        RECT 73.560 101.630 73.790 101.920 ;
        RECT 73.605 101.000 73.745 101.630 ;
        RECT 72.540 100.710 72.770 101.000 ;
        RECT 73.560 100.710 73.790 101.000 ;
        RECT 72.585 100.095 72.725 100.710 ;
        RECT 72.880 100.465 73.110 100.540 ;
        RECT 72.880 100.325 73.405 100.465 ;
        RECT 72.880 100.250 73.110 100.325 ;
        RECT 72.525 99.775 72.785 100.095 ;
        RECT 72.585 98.240 72.725 99.775 ;
        RECT 72.540 97.950 72.770 98.240 ;
        RECT 72.880 96.110 73.110 96.400 ;
        RECT 72.925 95.955 73.065 96.110 ;
        RECT 72.865 95.635 73.125 95.955 ;
        RECT 71.860 93.350 72.090 93.640 ;
        RECT 71.905 88.135 72.045 93.350 ;
        RECT 72.865 92.415 73.125 92.735 ;
        RECT 72.525 88.275 72.785 88.595 ;
        RECT 71.845 87.815 72.105 88.135 ;
        RECT 72.585 87.200 72.725 88.275 ;
        RECT 72.540 86.910 72.770 87.200 ;
        RECT 71.845 85.975 72.105 86.295 ;
        RECT 71.845 85.055 72.105 85.375 ;
        RECT 72.200 84.365 72.430 84.440 ;
        RECT 72.925 84.365 73.065 92.415 ;
        RECT 72.200 84.225 73.065 84.365 ;
        RECT 72.200 84.150 72.430 84.225 ;
        RECT 72.245 83.995 72.385 84.150 ;
        RECT 72.185 83.675 72.445 83.995 ;
        RECT 72.525 83.445 72.785 83.535 ;
        RECT 73.265 83.445 73.405 100.325 ;
        RECT 73.545 86.895 73.805 87.215 ;
        RECT 73.605 85.360 73.745 86.895 ;
        RECT 73.560 85.070 73.790 85.360 ;
        RECT 72.525 83.305 73.405 83.445 ;
        RECT 72.525 83.215 72.785 83.305 ;
        RECT 72.185 82.755 72.445 83.075 ;
        RECT 71.845 82.295 72.105 82.615 ;
        RECT 71.860 82.065 72.090 82.140 ;
        RECT 72.245 82.065 72.385 82.755 ;
        RECT 71.860 81.925 72.385 82.065 ;
        RECT 71.860 81.850 72.090 81.925 ;
        RECT 72.185 81.375 72.445 81.695 ;
        RECT 71.845 80.915 72.105 81.235 ;
        RECT 72.525 79.995 72.785 80.315 ;
        RECT 71.860 79.550 72.090 79.840 ;
        RECT 71.905 73.415 72.045 79.550 ;
        RECT 71.845 73.095 72.105 73.415 ;
        RECT 73.945 65.665 74.425 117.645 ;
        RECT 74.565 114.035 74.825 114.355 ;
        RECT 75.600 114.265 75.830 114.340 ;
        RECT 75.600 114.125 76.125 114.265 ;
        RECT 75.600 114.050 75.830 114.125 ;
        RECT 74.625 113.880 74.765 114.035 ;
        RECT 74.580 113.590 74.810 113.880 ;
        RECT 75.985 113.435 76.125 114.125 ;
        RECT 75.925 113.115 76.185 113.435 ;
        RECT 75.245 112.655 75.505 112.975 ;
        RECT 74.565 111.275 74.825 111.595 ;
        RECT 74.920 109.665 75.150 109.740 ;
        RECT 75.305 109.665 75.445 112.655 ;
        RECT 75.585 111.735 75.845 112.055 ;
        RECT 75.645 111.580 75.785 111.735 ;
        RECT 75.600 111.290 75.830 111.580 ;
        RECT 75.585 110.815 75.845 111.135 ;
        RECT 74.920 109.525 75.445 109.665 ;
        RECT 74.920 109.450 75.150 109.525 ;
        RECT 75.985 108.835 76.125 113.115 ;
        RECT 75.925 108.515 76.185 108.835 ;
        RECT 75.925 98.855 76.185 99.175 ;
        RECT 74.565 89.655 74.825 89.975 ;
        RECT 75.985 89.960 76.125 98.855 ;
        RECT 76.265 91.955 76.525 92.275 ;
        RECT 76.325 90.880 76.465 91.955 ;
        RECT 76.280 90.590 76.510 90.880 ;
        RECT 75.940 89.670 76.170 89.960 ;
        RECT 75.925 88.735 76.185 89.055 ;
        RECT 75.940 80.930 76.170 81.220 ;
        RECT 75.985 80.775 76.125 80.930 ;
        RECT 75.925 80.455 76.185 80.775 ;
        RECT 75.245 79.995 75.505 80.315 ;
        RECT 75.940 80.010 76.170 80.300 ;
        RECT 75.305 79.305 75.445 79.995 ;
        RECT 75.985 79.855 76.125 80.010 ;
        RECT 75.925 79.535 76.185 79.855 ;
        RECT 75.600 79.305 75.830 79.380 ;
        RECT 75.305 79.165 75.830 79.305 ;
        RECT 75.600 79.090 75.830 79.165 ;
        RECT 76.665 65.665 77.145 117.645 ;
        RECT 78.305 115.875 78.565 116.195 ;
        RECT 77.640 114.510 77.870 114.800 ;
        RECT 77.685 114.355 77.825 114.510 ;
        RECT 77.625 114.035 77.885 114.355 ;
        RECT 77.965 113.575 78.225 113.895 ;
        RECT 77.980 113.345 78.210 113.420 ;
        RECT 78.365 113.345 78.505 115.875 ;
        RECT 78.985 115.415 79.245 115.735 ;
        RECT 79.045 114.800 79.185 115.415 ;
        RECT 79.000 114.510 79.230 114.800 ;
        RECT 77.980 113.205 78.505 113.345 ;
        RECT 77.980 113.130 78.210 113.205 ;
        RECT 77.300 112.210 77.530 112.500 ;
        RECT 77.345 111.595 77.485 112.210 ;
        RECT 77.285 111.275 77.545 111.595 ;
        RECT 78.025 109.295 78.165 113.130 ;
        RECT 77.965 108.975 78.225 109.295 ;
        RECT 77.965 92.415 78.225 92.735 ;
        RECT 78.025 91.800 78.165 92.415 ;
        RECT 77.980 91.510 78.210 91.800 ;
        RECT 77.965 90.575 78.225 90.895 ;
        RECT 79.000 89.650 79.230 89.940 ;
        RECT 79.045 89.020 79.185 89.650 ;
        RECT 79.000 88.730 79.230 89.020 ;
        RECT 78.305 86.435 78.565 86.755 ;
        RECT 77.625 83.675 77.885 83.995 ;
        RECT 77.685 81.680 77.825 83.675 ;
        RECT 77.640 81.390 77.870 81.680 ;
        RECT 77.285 80.455 77.545 80.775 ;
        RECT 77.285 79.305 77.545 79.395 ;
        RECT 77.685 79.305 77.825 81.390 ;
        RECT 78.645 80.915 78.905 81.235 ;
        RECT 78.705 79.855 78.845 80.915 ;
        RECT 79.000 80.470 79.230 80.760 ;
        RECT 78.645 79.535 78.905 79.855 ;
        RECT 77.285 79.165 77.825 79.305 ;
        RECT 77.285 79.075 77.545 79.165 ;
        RECT 77.980 79.090 78.210 79.380 ;
        RECT 77.345 75.255 77.485 79.075 ;
        RECT 78.025 77.180 78.165 79.090 ;
        RECT 78.305 78.155 78.565 78.475 ;
        RECT 78.705 78.385 78.845 79.535 ;
        RECT 79.045 78.935 79.185 80.470 ;
        RECT 78.985 78.615 79.245 78.935 ;
        RECT 78.705 78.245 79.185 78.385 ;
        RECT 78.660 77.685 78.890 77.975 ;
        RECT 78.320 77.290 78.550 77.580 ;
        RECT 77.980 76.890 78.210 77.180 ;
        RECT 78.365 76.390 78.505 77.290 ;
        RECT 78.320 76.100 78.550 76.390 ;
        RECT 77.285 74.935 77.545 75.255 ;
        RECT 78.365 73.870 78.505 76.100 ;
        RECT 78.705 75.875 78.845 77.685 ;
        RECT 79.045 77.095 79.185 78.245 ;
        RECT 78.985 76.775 79.245 77.095 ;
        RECT 78.660 75.585 78.890 75.875 ;
        RECT 78.705 74.305 78.845 75.585 ;
        RECT 78.660 74.015 78.890 74.305 ;
        RECT 78.320 73.580 78.550 73.870 ;
        RECT 79.045 71.560 79.185 76.775 ;
        RECT 79.000 71.270 79.230 71.560 ;
        RECT 79.385 65.665 79.865 117.645 ;
        RECT 81.025 115.875 81.285 116.195 ;
        RECT 81.720 115.185 81.950 115.260 ;
        RECT 81.425 115.045 81.950 115.185 ;
        RECT 81.040 114.510 81.270 114.800 ;
        RECT 81.085 113.895 81.225 114.510 ;
        RECT 81.025 113.575 81.285 113.895 ;
        RECT 81.040 113.130 81.270 113.420 ;
        RECT 81.085 112.975 81.225 113.130 ;
        RECT 80.360 112.645 80.590 112.935 ;
        RECT 81.025 112.655 81.285 112.975 ;
        RECT 80.405 110.835 80.545 112.645 ;
        RECT 80.700 112.250 80.930 112.540 ;
        RECT 80.745 111.350 80.885 112.250 ;
        RECT 81.425 112.085 81.565 115.045 ;
        RECT 81.720 114.970 81.950 115.045 ;
        RECT 81.720 113.590 81.950 113.880 ;
        RECT 81.765 112.515 81.905 113.590 ;
        RECT 81.705 112.195 81.965 112.515 ;
        RECT 81.380 111.795 81.610 112.085 ;
        RECT 80.700 111.060 80.930 111.350 ;
        RECT 80.360 110.545 80.590 110.835 ;
        RECT 80.405 109.265 80.545 110.545 ;
        RECT 80.360 108.975 80.590 109.265 ;
        RECT 80.745 108.830 80.885 111.060 ;
        RECT 80.700 108.540 80.930 108.830 ;
        RECT 80.360 106.230 80.590 106.520 ;
        RECT 80.005 102.765 80.265 102.855 ;
        RECT 80.405 102.765 80.545 106.230 ;
        RECT 81.720 103.930 81.950 104.220 ;
        RECT 81.025 103.455 81.285 103.775 ;
        RECT 81.085 103.300 81.225 103.455 ;
        RECT 81.040 103.225 81.270 103.300 ;
        RECT 81.040 103.085 81.565 103.225 ;
        RECT 81.040 103.010 81.270 103.085 ;
        RECT 80.005 102.625 80.545 102.765 ;
        RECT 80.005 102.535 80.265 102.625 ;
        RECT 81.040 102.305 81.270 102.380 ;
        RECT 80.745 102.165 81.270 102.305 ;
        RECT 80.020 101.630 80.250 101.920 ;
        RECT 80.065 101.000 80.205 101.630 ;
        RECT 80.020 100.710 80.250 101.000 ;
        RECT 80.745 100.005 80.885 102.165 ;
        RECT 81.040 102.090 81.270 102.165 ;
        RECT 81.040 101.385 81.270 101.460 ;
        RECT 81.425 101.385 81.565 103.085 ;
        RECT 81.040 101.245 81.565 101.385 ;
        RECT 81.040 101.170 81.270 101.245 ;
        RECT 81.040 100.710 81.270 101.000 ;
        RECT 81.085 100.095 81.225 100.710 ;
        RECT 81.025 100.005 81.285 100.095 ;
        RECT 80.745 99.865 81.285 100.005 ;
        RECT 81.025 99.775 81.285 99.865 ;
        RECT 81.085 98.240 81.225 99.775 ;
        RECT 81.765 99.175 81.905 103.930 ;
        RECT 81.705 98.855 81.965 99.175 ;
        RECT 81.040 97.950 81.270 98.240 ;
        RECT 80.700 96.110 80.930 96.400 ;
        RECT 80.020 94.270 80.250 94.560 ;
        RECT 80.065 93.195 80.205 94.270 ;
        RECT 80.005 92.875 80.265 93.195 ;
        RECT 80.745 92.735 80.885 96.110 ;
        RECT 81.705 95.175 81.965 95.495 ;
        RECT 81.720 94.270 81.950 94.560 ;
        RECT 81.765 94.115 81.905 94.270 ;
        RECT 81.705 93.795 81.965 94.115 ;
        RECT 81.365 93.335 81.625 93.655 ;
        RECT 80.685 92.415 80.945 92.735 ;
        RECT 81.705 91.495 81.965 91.815 ;
        RECT 81.765 90.895 81.905 91.495 ;
        RECT 81.705 90.575 81.965 90.895 ;
        RECT 80.700 88.280 80.930 88.570 ;
        RECT 80.360 87.845 80.590 88.135 ;
        RECT 80.405 86.565 80.545 87.845 ;
        RECT 80.360 86.275 80.590 86.565 ;
        RECT 80.405 84.465 80.545 86.275 ;
        RECT 80.745 86.050 80.885 88.280 ;
        RECT 81.025 86.435 81.285 86.755 ;
        RECT 80.700 85.760 80.930 86.050 ;
        RECT 80.745 84.860 80.885 85.760 ;
        RECT 81.085 85.315 81.225 86.435 ;
        RECT 81.040 85.025 81.270 85.315 ;
        RECT 80.700 84.570 80.930 84.860 ;
        RECT 80.360 84.175 80.590 84.465 ;
        RECT 80.700 83.690 80.930 83.980 ;
        RECT 80.745 82.155 80.885 83.690 ;
        RECT 80.685 81.835 80.945 82.155 ;
        RECT 80.005 80.455 80.265 80.775 ;
        RECT 80.065 80.300 80.205 80.455 ;
        RECT 80.020 80.010 80.250 80.300 ;
        RECT 80.005 78.615 80.265 78.935 ;
        RECT 80.065 78.000 80.205 78.615 ;
        RECT 80.345 78.385 80.605 78.475 ;
        RECT 80.745 78.385 80.885 81.835 ;
        RECT 81.365 80.915 81.625 81.235 ;
        RECT 81.365 80.225 81.625 80.315 ;
        RECT 81.085 80.085 81.625 80.225 ;
        RECT 81.085 78.460 81.225 80.085 ;
        RECT 81.365 79.995 81.625 80.085 ;
        RECT 81.720 79.090 81.950 79.380 ;
        RECT 80.345 78.245 80.885 78.385 ;
        RECT 80.345 78.155 80.605 78.245 ;
        RECT 81.040 78.170 81.270 78.460 ;
        RECT 80.020 77.710 80.250 78.000 ;
        RECT 81.025 76.775 81.285 77.095 ;
        RECT 81.765 73.875 81.905 79.090 ;
        RECT 81.705 73.555 81.965 73.875 ;
        RECT 82.105 65.665 82.585 117.645 ;
        RECT 83.420 113.590 83.650 113.880 ;
        RECT 83.465 113.435 83.605 113.590 ;
        RECT 83.405 113.115 83.665 113.435 ;
        RECT 84.100 113.105 84.330 113.395 ;
        RECT 83.760 112.710 83.990 113.000 ;
        RECT 83.080 112.515 83.310 112.545 ;
        RECT 83.065 112.195 83.325 112.515 ;
        RECT 83.805 111.810 83.945 112.710 ;
        RECT 83.760 111.520 83.990 111.810 ;
        RECT 83.805 109.290 83.945 111.520 ;
        RECT 84.145 111.295 84.285 113.105 ;
        RECT 84.100 111.005 84.330 111.295 ;
        RECT 84.145 109.725 84.285 111.005 ;
        RECT 84.100 109.435 84.330 109.725 ;
        RECT 83.760 109.000 83.990 109.290 ;
        RECT 84.440 106.690 84.670 106.980 ;
        RECT 84.485 106.535 84.625 106.690 ;
        RECT 84.425 106.215 84.685 106.535 ;
        RECT 83.745 103.455 84.005 103.775 ;
        RECT 83.420 103.010 83.650 103.300 ;
        RECT 83.465 102.855 83.605 103.010 ;
        RECT 83.405 102.535 83.665 102.855 ;
        RECT 83.805 102.380 83.945 103.455 ;
        RECT 83.760 102.090 83.990 102.380 ;
        RECT 83.420 101.170 83.650 101.460 ;
        RECT 84.100 101.170 84.330 101.460 ;
        RECT 83.465 100.095 83.605 101.170 ;
        RECT 84.145 100.095 84.285 101.170 ;
        RECT 83.405 99.775 83.665 100.095 ;
        RECT 84.085 99.775 84.345 100.095 ;
        RECT 84.440 97.950 84.670 98.240 ;
        RECT 84.485 96.875 84.625 97.950 ;
        RECT 83.405 96.555 83.665 96.875 ;
        RECT 84.425 96.555 84.685 96.875 ;
        RECT 83.420 96.325 83.650 96.400 ;
        RECT 83.125 96.185 83.650 96.325 ;
        RECT 82.740 94.730 82.970 95.020 ;
        RECT 82.785 89.975 82.925 94.730 ;
        RECT 83.125 92.275 83.265 96.185 ;
        RECT 83.420 96.110 83.650 96.185 ;
        RECT 83.405 95.635 83.665 95.955 ;
        RECT 83.760 94.270 83.990 94.560 ;
        RECT 83.405 92.415 83.665 92.735 ;
        RECT 83.805 92.275 83.945 94.270 ;
        RECT 83.065 91.955 83.325 92.275 ;
        RECT 83.745 91.955 84.005 92.275 ;
        RECT 83.420 90.590 83.650 90.880 ;
        RECT 82.725 89.655 82.985 89.975 ;
        RECT 83.080 82.065 83.310 82.140 ;
        RECT 82.785 81.925 83.310 82.065 ;
        RECT 82.785 80.315 82.925 81.925 ;
        RECT 83.080 81.850 83.310 81.925 ;
        RECT 83.465 81.680 83.605 90.590 ;
        RECT 84.440 90.570 84.670 90.860 ;
        RECT 84.485 89.940 84.625 90.570 ;
        RECT 84.440 89.650 84.670 89.940 ;
        RECT 83.745 87.815 84.005 88.135 ;
        RECT 83.420 81.390 83.650 81.680 ;
        RECT 83.465 81.235 83.605 81.390 ;
        RECT 83.405 80.915 83.665 81.235 ;
        RECT 83.405 80.685 83.665 80.775 ;
        RECT 83.125 80.545 83.665 80.685 ;
        RECT 82.725 79.995 82.985 80.315 ;
        RECT 82.740 71.025 82.970 71.100 ;
        RECT 83.125 71.025 83.265 80.545 ;
        RECT 83.405 80.455 83.665 80.545 ;
        RECT 84.440 79.550 84.670 79.840 ;
        RECT 83.405 78.155 83.665 78.475 ;
        RECT 83.465 78.000 83.605 78.155 ;
        RECT 84.485 78.015 84.625 79.550 ;
        RECT 83.420 77.710 83.650 78.000 ;
        RECT 84.425 77.695 84.685 78.015 ;
        RECT 84.100 77.225 84.330 77.515 ;
        RECT 83.760 76.830 83.990 77.120 ;
        RECT 83.420 76.635 83.650 76.665 ;
        RECT 83.405 76.315 83.665 76.635 ;
        RECT 83.805 75.930 83.945 76.830 ;
        RECT 83.760 75.640 83.990 75.930 ;
        RECT 83.805 73.410 83.945 75.640 ;
        RECT 84.145 75.415 84.285 77.225 ;
        RECT 84.100 75.125 84.330 75.415 ;
        RECT 84.145 73.845 84.285 75.125 ;
        RECT 84.100 73.555 84.330 73.845 ;
        RECT 83.760 73.120 83.990 73.410 ;
        RECT 82.740 70.885 83.265 71.025 ;
        RECT 82.740 70.810 82.970 70.885 ;
        RECT 84.825 65.665 85.305 117.645 ;
        RECT 86.805 106.215 87.065 106.535 ;
        RECT 86.125 105.755 86.385 106.075 ;
        RECT 85.460 104.850 85.690 105.140 ;
        RECT 85.505 103.775 85.645 104.850 ;
        RECT 86.465 104.835 86.725 105.155 ;
        RECT 87.145 103.915 87.405 104.235 ;
        RECT 85.445 103.455 85.705 103.775 ;
        RECT 85.800 103.225 86.030 103.300 ;
        RECT 85.505 103.085 86.030 103.225 ;
        RECT 85.505 96.325 85.645 103.085 ;
        RECT 85.800 103.010 86.030 103.085 ;
        RECT 86.480 102.305 86.710 102.380 ;
        RECT 86.185 102.165 86.710 102.305 ;
        RECT 86.185 100.095 86.325 102.165 ;
        RECT 86.480 102.090 86.710 102.165 ;
        RECT 87.160 101.845 87.390 101.920 ;
        RECT 86.525 101.705 87.390 101.845 ;
        RECT 86.125 99.775 86.385 100.095 ;
        RECT 86.525 99.175 86.665 101.705 ;
        RECT 87.160 101.630 87.390 101.705 ;
        RECT 87.160 101.170 87.390 101.460 ;
        RECT 86.820 100.250 87.050 100.540 ;
        RECT 86.865 100.095 87.005 100.250 ;
        RECT 86.805 99.775 87.065 100.095 ;
        RECT 87.205 99.545 87.345 101.170 ;
        RECT 86.865 99.405 87.345 99.545 ;
        RECT 86.465 98.855 86.725 99.175 ;
        RECT 86.480 97.245 86.710 97.320 ;
        RECT 86.865 97.245 87.005 99.405 ;
        RECT 87.145 98.855 87.405 99.175 ;
        RECT 86.480 97.105 87.005 97.245 ;
        RECT 86.480 97.030 86.710 97.105 ;
        RECT 86.465 96.555 86.725 96.875 ;
        RECT 86.140 96.325 86.370 96.400 ;
        RECT 85.505 96.185 86.370 96.325 ;
        RECT 86.140 96.110 86.370 96.185 ;
        RECT 85.460 95.650 85.690 95.940 ;
        RECT 86.865 95.865 87.005 97.105 ;
        RECT 86.185 95.725 87.005 95.865 ;
        RECT 85.505 95.495 85.645 95.650 ;
        RECT 85.445 95.175 85.705 95.495 ;
        RECT 85.785 80.915 86.045 81.235 ;
        RECT 85.845 78.920 85.985 80.915 ;
        RECT 86.185 80.775 86.325 95.725 ;
        RECT 86.480 95.190 86.710 95.480 ;
        RECT 86.525 95.035 86.665 95.190 ;
        RECT 86.465 94.715 86.725 95.035 ;
        RECT 87.160 94.270 87.390 94.560 ;
        RECT 86.805 93.335 87.065 93.655 ;
        RECT 86.465 91.035 86.725 91.355 ;
        RECT 86.125 80.455 86.385 80.775 ;
        RECT 86.185 79.765 86.325 80.455 ;
        RECT 86.480 80.225 86.710 80.300 ;
        RECT 86.865 80.225 87.005 93.335 ;
        RECT 87.205 90.435 87.345 94.270 ;
        RECT 87.145 90.115 87.405 90.435 ;
        RECT 87.145 88.275 87.405 88.595 ;
        RECT 87.205 84.900 87.345 88.275 ;
        RECT 87.160 84.610 87.390 84.900 ;
        RECT 87.145 81.375 87.405 81.695 ;
        RECT 87.160 80.470 87.390 80.760 ;
        RECT 87.205 80.315 87.345 80.470 ;
        RECT 86.480 80.085 87.005 80.225 ;
        RECT 86.480 80.010 86.710 80.085 ;
        RECT 86.480 79.765 86.710 79.840 ;
        RECT 86.185 79.625 86.710 79.765 ;
        RECT 86.480 79.550 86.710 79.625 ;
        RECT 85.800 78.630 86.030 78.920 ;
        RECT 86.865 78.845 87.005 80.085 ;
        RECT 87.145 79.995 87.405 80.315 ;
        RECT 87.145 79.535 87.405 79.855 ;
        RECT 86.525 78.705 87.005 78.845 ;
        RECT 85.460 77.465 85.690 77.540 ;
        RECT 85.460 77.325 85.985 77.465 ;
        RECT 85.460 77.250 85.690 77.325 ;
        RECT 85.445 76.315 85.705 76.635 ;
        RECT 85.845 72.940 85.985 77.325 ;
        RECT 86.525 74.705 86.665 78.705 ;
        RECT 86.820 78.385 87.050 78.460 ;
        RECT 87.205 78.385 87.345 79.535 ;
        RECT 86.820 78.245 87.345 78.385 ;
        RECT 86.820 78.170 87.050 78.245 ;
        RECT 86.805 77.695 87.065 78.015 ;
        RECT 86.865 77.540 87.005 77.695 ;
        RECT 86.820 77.250 87.050 77.540 ;
        RECT 86.805 76.315 87.065 76.635 ;
        RECT 86.865 75.700 87.005 76.315 ;
        RECT 86.820 75.410 87.050 75.700 ;
        RECT 86.805 74.705 87.065 74.795 ;
        RECT 86.525 74.565 87.065 74.705 ;
        RECT 86.805 74.475 87.065 74.565 ;
        RECT 86.465 73.555 86.725 73.875 ;
        RECT 86.525 73.400 86.665 73.555 ;
        RECT 86.480 73.110 86.710 73.400 ;
        RECT 85.800 72.650 86.030 72.940 ;
        RECT 87.545 65.665 88.025 117.645 ;
        RECT 88.860 115.890 89.090 116.180 ;
        RECT 88.905 115.735 89.045 115.890 ;
        RECT 88.845 115.415 89.105 115.735 ;
        RECT 88.180 115.185 88.410 115.260 ;
        RECT 88.180 115.045 88.705 115.185 ;
        RECT 88.180 114.970 88.410 115.045 ;
        RECT 88.565 113.575 88.705 115.045 ;
        RECT 88.520 113.285 88.750 113.575 ;
        RECT 88.905 109.295 89.045 115.415 ;
        RECT 89.185 114.495 89.445 114.815 ;
        RECT 89.540 114.025 89.770 114.315 ;
        RECT 89.200 113.630 89.430 113.920 ;
        RECT 89.245 112.730 89.385 113.630 ;
        RECT 89.200 112.440 89.430 112.730 ;
        RECT 89.245 110.210 89.385 112.440 ;
        RECT 89.585 112.215 89.725 114.025 ;
        RECT 89.540 111.925 89.770 112.215 ;
        RECT 89.585 110.645 89.725 111.925 ;
        RECT 89.540 110.355 89.770 110.645 ;
        RECT 89.200 109.920 89.430 110.210 ;
        RECT 88.845 108.975 89.105 109.295 ;
        RECT 88.180 107.610 88.410 107.900 ;
        RECT 88.225 105.155 88.365 107.610 ;
        RECT 88.505 105.755 88.765 106.075 ;
        RECT 88.165 104.835 88.425 105.155 ;
        RECT 88.165 103.455 88.425 103.775 ;
        RECT 88.225 101.475 88.365 103.455 ;
        RECT 88.165 101.155 88.425 101.475 ;
        RECT 88.225 99.635 88.365 101.155 ;
        RECT 88.565 100.925 88.705 105.755 ;
        RECT 88.845 104.835 89.105 105.155 ;
        RECT 88.905 103.300 89.045 104.835 ;
        RECT 88.860 103.225 89.090 103.300 ;
        RECT 88.860 103.085 89.385 103.225 ;
        RECT 88.860 103.010 89.090 103.085 ;
        RECT 88.845 102.535 89.105 102.855 ;
        RECT 88.845 101.155 89.105 101.475 ;
        RECT 89.245 101.385 89.385 103.085 ;
        RECT 89.865 102.535 90.125 102.855 ;
        RECT 89.245 101.245 89.725 101.385 ;
        RECT 88.565 100.785 89.385 100.925 ;
        RECT 88.565 100.080 88.705 100.785 ;
        RECT 88.860 100.250 89.090 100.540 ;
        RECT 88.520 99.790 88.750 100.080 ;
        RECT 88.165 99.545 88.425 99.635 ;
        RECT 88.165 99.405 88.705 99.545 ;
        RECT 88.165 99.315 88.425 99.405 ;
        RECT 88.165 98.395 88.425 98.715 ;
        RECT 88.225 94.115 88.365 98.395 ;
        RECT 88.565 96.000 88.705 99.405 ;
        RECT 88.905 99.160 89.045 100.250 ;
        RECT 88.860 98.870 89.090 99.160 ;
        RECT 88.905 98.715 89.045 98.870 ;
        RECT 88.845 98.395 89.105 98.715 ;
        RECT 88.845 97.935 89.105 98.255 ;
        RECT 88.845 97.015 89.105 97.335 ;
        RECT 88.885 96.860 89.025 97.015 ;
        RECT 88.860 96.570 89.090 96.860 ;
        RECT 88.860 96.110 89.090 96.400 ;
        RECT 88.520 95.710 88.750 96.000 ;
        RECT 88.905 94.945 89.045 96.110 ;
        RECT 89.245 95.480 89.385 100.785 ;
        RECT 89.200 95.190 89.430 95.480 ;
        RECT 88.905 94.805 89.385 94.945 ;
        RECT 88.860 94.270 89.090 94.560 ;
        RECT 88.165 93.795 88.425 94.115 ;
        RECT 88.905 93.105 89.045 94.270 ;
        RECT 89.245 93.655 89.385 94.805 ;
        RECT 89.185 93.335 89.445 93.655 ;
        RECT 89.585 93.105 89.725 101.245 ;
        RECT 89.925 95.940 90.065 102.535 ;
        RECT 89.880 95.650 90.110 95.940 ;
        RECT 89.865 93.795 90.125 94.115 ;
        RECT 89.925 93.640 90.065 93.795 ;
        RECT 89.880 93.350 90.110 93.640 ;
        RECT 89.925 93.195 90.065 93.350 ;
        RECT 88.905 92.965 89.725 93.105 ;
        RECT 89.865 92.875 90.125 93.195 ;
        RECT 88.845 92.415 89.105 92.735 ;
        RECT 88.905 91.340 89.045 92.415 ;
        RECT 89.865 91.955 90.125 92.275 ;
        RECT 89.925 91.340 90.065 91.955 ;
        RECT 88.860 91.050 89.090 91.340 ;
        RECT 89.880 91.050 90.110 91.340 ;
        RECT 88.845 90.115 89.105 90.435 ;
        RECT 88.860 89.670 89.090 89.960 ;
        RECT 88.905 88.135 89.045 89.670 ;
        RECT 89.540 88.750 89.770 89.040 ;
        RECT 88.845 87.815 89.105 88.135 ;
        RECT 89.585 85.375 89.725 88.750 ;
        RECT 89.525 85.285 89.785 85.375 ;
        RECT 88.565 85.145 89.785 85.285 ;
        RECT 88.565 81.680 88.705 85.145 ;
        RECT 89.525 85.055 89.785 85.145 ;
        RECT 88.520 81.390 88.750 81.680 ;
        RECT 88.180 80.470 88.410 80.760 ;
        RECT 88.225 76.635 88.365 80.470 ;
        RECT 88.565 79.855 88.705 81.390 ;
        RECT 89.185 81.375 89.445 81.695 ;
        RECT 88.505 79.535 88.765 79.855 ;
        RECT 88.860 79.305 89.090 79.380 ;
        RECT 88.565 79.165 89.090 79.305 ;
        RECT 88.165 76.315 88.425 76.635 ;
        RECT 88.565 75.855 88.705 79.165 ;
        RECT 88.860 79.090 89.090 79.165 ;
        RECT 89.245 78.935 89.385 81.375 ;
        RECT 89.880 80.470 90.110 80.760 ;
        RECT 89.185 78.845 89.445 78.935 ;
        RECT 88.905 78.705 89.445 78.845 ;
        RECT 88.905 77.540 89.045 78.705 ;
        RECT 89.185 78.615 89.445 78.705 ;
        RECT 89.185 77.695 89.445 78.015 ;
        RECT 89.925 78.000 90.065 80.470 ;
        RECT 89.880 77.710 90.110 78.000 ;
        RECT 88.860 77.250 89.090 77.540 ;
        RECT 89.245 77.080 89.385 77.695 ;
        RECT 89.200 76.790 89.430 77.080 ;
        RECT 89.540 76.305 89.770 76.595 ;
        RECT 89.200 75.910 89.430 76.200 ;
        RECT 88.520 75.565 88.750 75.855 ;
        RECT 89.245 75.010 89.385 75.910 ;
        RECT 88.165 74.475 88.425 74.795 ;
        RECT 89.200 74.720 89.430 75.010 ;
        RECT 88.225 70.180 88.365 74.475 ;
        RECT 89.245 72.490 89.385 74.720 ;
        RECT 89.585 74.495 89.725 76.305 ;
        RECT 89.540 74.205 89.770 74.495 ;
        RECT 89.585 72.925 89.725 74.205 ;
        RECT 89.540 72.635 89.770 72.925 ;
        RECT 89.200 72.200 89.430 72.490 ;
        RECT 88.180 69.890 88.410 70.180 ;
        RECT 90.265 65.665 90.745 117.645 ;
        RECT 91.920 115.890 92.150 116.180 ;
        RECT 91.965 115.735 92.105 115.890 ;
        RECT 91.905 115.415 92.165 115.735 ;
        RECT 91.240 115.185 91.470 115.260 ;
        RECT 91.240 115.045 91.765 115.185 ;
        RECT 91.240 114.970 91.470 115.045 ;
        RECT 91.240 114.025 91.470 114.315 ;
        RECT 91.625 114.265 91.765 115.045 ;
        RECT 91.905 114.725 92.165 114.815 ;
        RECT 91.905 114.585 92.445 114.725 ;
        RECT 91.905 114.495 92.165 114.585 ;
        RECT 91.625 114.125 92.105 114.265 ;
        RECT 91.285 112.215 91.425 114.025 ;
        RECT 91.580 113.630 91.810 113.920 ;
        RECT 91.625 112.730 91.765 113.630 ;
        RECT 91.965 113.520 92.105 114.125 ;
        RECT 91.920 113.230 92.150 113.520 ;
        RECT 92.305 113.345 92.445 114.585 ;
        RECT 92.585 113.345 92.845 113.435 ;
        RECT 92.305 113.205 92.845 113.345 ;
        RECT 92.585 113.115 92.845 113.205 ;
        RECT 91.580 112.440 91.810 112.730 ;
        RECT 91.240 111.925 91.470 112.215 ;
        RECT 91.285 110.645 91.425 111.925 ;
        RECT 91.240 110.355 91.470 110.645 ;
        RECT 91.625 110.210 91.765 112.440 ;
        RECT 91.580 109.920 91.810 110.210 ;
        RECT 90.900 107.610 91.130 107.900 ;
        RECT 90.945 106.075 91.085 107.610 ;
        RECT 91.905 106.215 92.165 106.535 ;
        RECT 90.885 105.755 91.145 106.075 ;
        RECT 91.580 104.390 91.810 104.680 ;
        RECT 91.625 104.235 91.765 104.390 ;
        RECT 90.900 103.930 91.130 104.220 ;
        RECT 90.945 103.775 91.085 103.930 ;
        RECT 91.565 103.915 91.825 104.235 ;
        RECT 90.885 103.455 91.145 103.775 ;
        RECT 91.965 102.370 92.105 106.215 ;
        RECT 91.920 102.080 92.150 102.370 ;
        RECT 92.600 102.090 92.830 102.380 ;
        RECT 91.240 101.170 91.470 101.460 ;
        RECT 90.885 99.315 91.145 99.635 ;
        RECT 90.945 98.240 91.085 99.315 ;
        RECT 90.900 97.950 91.130 98.240 ;
        RECT 90.885 97.475 91.145 97.795 ;
        RECT 90.945 94.115 91.085 97.475 ;
        RECT 90.885 93.795 91.145 94.115 ;
        RECT 90.885 93.335 91.145 93.655 ;
        RECT 90.885 92.415 91.145 92.735 ;
        RECT 90.900 88.770 91.130 89.060 ;
        RECT 90.945 88.140 91.085 88.770 ;
        RECT 91.285 88.505 91.425 101.170 ;
        RECT 91.905 98.855 92.165 99.175 ;
        RECT 91.965 98.240 92.105 98.855 ;
        RECT 92.645 98.255 92.785 102.090 ;
        RECT 91.920 97.950 92.150 98.240 ;
        RECT 92.585 97.935 92.845 98.255 ;
        RECT 91.580 97.030 91.810 97.320 ;
        RECT 91.625 95.955 91.765 97.030 ;
        RECT 91.905 96.555 92.165 96.875 ;
        RECT 91.565 95.635 91.825 95.955 ;
        RECT 92.600 95.650 92.830 95.940 ;
        RECT 92.260 94.945 92.490 95.020 ;
        RECT 92.645 94.945 92.785 95.650 ;
        RECT 92.260 94.805 92.785 94.945 ;
        RECT 92.260 94.730 92.490 94.805 ;
        RECT 91.580 93.810 91.810 94.100 ;
        RECT 91.625 93.195 91.765 93.810 ;
        RECT 91.920 93.350 92.150 93.640 ;
        RECT 91.565 92.875 91.825 93.195 ;
        RECT 91.965 91.340 92.105 93.350 ;
        RECT 91.920 91.050 92.150 91.340 ;
        RECT 91.580 88.505 91.810 88.580 ;
        RECT 91.285 88.365 91.810 88.505 ;
        RECT 91.580 88.290 91.810 88.365 ;
        RECT 90.900 87.850 91.130 88.140 ;
        RECT 91.225 87.355 91.485 87.675 ;
        RECT 90.900 84.150 91.130 84.440 ;
        RECT 90.945 82.155 91.085 84.150 ;
        RECT 90.885 81.835 91.145 82.155 ;
        RECT 90.900 81.605 91.130 81.680 ;
        RECT 91.285 81.605 91.425 87.355 ;
        RECT 91.920 86.910 92.150 87.200 ;
        RECT 91.965 82.525 92.105 86.910 ;
        RECT 92.245 85.055 92.505 85.375 ;
        RECT 92.305 83.075 92.445 85.055 ;
        RECT 92.585 84.135 92.845 84.455 ;
        RECT 92.585 83.215 92.845 83.535 ;
        RECT 92.245 82.985 92.505 83.075 ;
        RECT 92.245 82.845 92.785 82.985 ;
        RECT 92.245 82.755 92.505 82.845 ;
        RECT 92.245 82.525 92.505 82.615 ;
        RECT 91.965 82.385 92.505 82.525 ;
        RECT 92.245 82.295 92.505 82.385 ;
        RECT 90.900 81.465 91.425 81.605 ;
        RECT 90.900 81.390 91.130 81.465 ;
        RECT 92.245 81.375 92.505 81.695 ;
        RECT 92.645 81.145 92.785 82.845 ;
        RECT 92.305 81.005 92.785 81.145 ;
        RECT 92.305 79.380 92.445 81.005 ;
        RECT 92.585 80.455 92.845 80.775 ;
        RECT 92.260 79.090 92.490 79.380 ;
        RECT 90.885 78.155 91.145 78.475 ;
        RECT 92.260 78.170 92.490 78.460 ;
        RECT 92.305 75.715 92.445 78.170 ;
        RECT 92.585 77.235 92.845 77.555 ;
        RECT 92.245 75.395 92.505 75.715 ;
        RECT 92.985 65.665 93.465 117.645 ;
        RECT 94.965 113.115 95.225 113.435 ;
        RECT 94.285 103.915 94.545 104.235 ;
        RECT 94.345 103.300 94.485 103.915 ;
        RECT 94.300 103.010 94.530 103.300 ;
        RECT 94.625 102.535 94.885 102.855 ;
        RECT 94.640 100.250 94.870 100.540 ;
        RECT 93.605 99.315 93.865 99.635 ;
        RECT 94.285 99.315 94.545 99.635 ;
        RECT 94.300 97.705 94.530 97.780 ;
        RECT 93.665 97.565 94.530 97.705 ;
        RECT 93.665 94.575 93.805 97.565 ;
        RECT 94.300 97.490 94.530 97.565 ;
        RECT 94.685 95.495 94.825 100.250 ;
        RECT 94.625 95.175 94.885 95.495 ;
        RECT 95.025 94.945 95.165 113.115 ;
        RECT 95.305 103.455 95.565 103.775 ;
        RECT 95.365 102.840 95.505 103.455 ;
        RECT 95.320 102.550 95.550 102.840 ;
        RECT 95.320 101.170 95.550 101.460 ;
        RECT 95.365 99.635 95.505 101.170 ;
        RECT 95.305 99.315 95.565 99.635 ;
        RECT 95.320 94.945 95.550 95.020 ;
        RECT 95.025 94.805 95.550 94.945 ;
        RECT 95.320 94.730 95.550 94.805 ;
        RECT 93.605 94.255 93.865 94.575 ;
        RECT 93.665 87.675 93.805 94.255 ;
        RECT 95.365 94.115 95.505 94.730 ;
        RECT 95.305 93.795 95.565 94.115 ;
        RECT 93.945 88.275 94.205 88.595 ;
        RECT 93.605 87.355 93.865 87.675 ;
        RECT 94.640 85.060 94.870 85.350 ;
        RECT 93.945 83.215 94.205 83.535 ;
        RECT 94.005 82.095 94.145 83.215 ;
        RECT 94.685 82.830 94.825 85.060 ;
        RECT 94.980 84.625 95.210 84.915 ;
        RECT 95.025 83.345 95.165 84.625 ;
        RECT 94.980 83.055 95.210 83.345 ;
        RECT 94.640 82.540 94.870 82.830 ;
        RECT 93.960 81.805 94.190 82.095 ;
        RECT 94.685 81.640 94.825 82.540 ;
        RECT 94.640 81.350 94.870 81.640 ;
        RECT 95.025 81.245 95.165 83.055 ;
        RECT 95.305 82.295 95.565 82.615 ;
        RECT 94.285 80.915 94.545 81.235 ;
        RECT 94.980 80.955 95.210 81.245 ;
        RECT 94.345 80.760 94.485 80.915 ;
        RECT 94.300 80.470 94.530 80.760 ;
        RECT 94.345 78.015 94.485 80.470 ;
        RECT 94.285 77.695 94.545 78.015 ;
        RECT 93.945 77.235 94.205 77.555 ;
        RECT 94.005 76.775 94.145 77.235 ;
        RECT 94.980 77.225 95.210 77.515 ;
        RECT 94.640 76.830 94.870 77.120 ;
        RECT 93.960 76.485 94.190 76.775 ;
        RECT 94.685 75.930 94.825 76.830 ;
        RECT 94.640 75.640 94.870 75.930 ;
        RECT 94.685 73.410 94.825 75.640 ;
        RECT 95.025 75.415 95.165 77.225 ;
        RECT 94.980 75.125 95.210 75.415 ;
        RECT 95.025 73.845 95.165 75.125 ;
        RECT 94.980 73.555 95.210 73.845 ;
        RECT 94.640 73.120 94.870 73.410 ;
        RECT 95.365 71.100 95.505 82.295 ;
        RECT 95.320 70.810 95.550 71.100 ;
        RECT 95.705 65.665 96.185 117.645 ;
        RECT 97.345 115.875 97.605 116.195 ;
        RECT 96.325 114.495 96.585 114.815 ;
        RECT 97.405 114.800 97.545 115.875 ;
        RECT 97.360 114.510 97.590 114.800 ;
        RECT 97.005 114.035 97.265 114.355 ;
        RECT 97.405 113.895 97.545 114.510 ;
        RECT 97.345 113.575 97.605 113.895 ;
        RECT 97.360 113.130 97.590 113.420 ;
        RECT 96.340 112.210 96.570 112.500 ;
        RECT 96.385 111.135 96.525 112.210 ;
        RECT 96.325 110.815 96.585 111.135 ;
        RECT 97.405 110.660 97.545 113.130 ;
        RECT 98.025 111.275 98.285 111.595 ;
        RECT 97.360 110.370 97.590 110.660 ;
        RECT 97.405 108.835 97.545 110.370 ;
        RECT 97.345 108.515 97.605 108.835 ;
        RECT 97.005 104.375 97.265 104.695 ;
        RECT 97.065 103.775 97.205 104.375 ;
        RECT 97.345 103.915 97.605 104.235 ;
        RECT 97.005 103.455 97.265 103.775 ;
        RECT 97.405 102.840 97.545 103.915 ;
        RECT 97.685 102.995 97.945 103.315 ;
        RECT 97.360 102.550 97.590 102.840 ;
        RECT 96.680 101.170 96.910 101.460 ;
        RECT 96.340 100.250 96.570 100.540 ;
        RECT 96.385 99.620 96.525 100.250 ;
        RECT 96.340 99.330 96.570 99.620 ;
        RECT 96.725 95.495 96.865 101.170 ;
        RECT 97.745 101.000 97.885 102.995 ;
        RECT 97.700 100.710 97.930 101.000 ;
        RECT 97.360 99.605 97.590 99.620 ;
        RECT 97.315 99.345 97.635 99.605 ;
        RECT 97.360 99.330 97.590 99.345 ;
        RECT 97.005 98.855 97.265 99.175 ;
        RECT 97.405 96.860 97.545 99.330 ;
        RECT 97.360 96.570 97.590 96.860 ;
        RECT 96.665 95.175 96.925 95.495 ;
        RECT 97.005 94.945 97.265 95.035 ;
        RECT 97.005 94.805 97.545 94.945 ;
        RECT 97.005 94.715 97.265 94.805 ;
        RECT 97.005 93.335 97.265 93.655 ;
        RECT 97.065 91.340 97.205 93.335 ;
        RECT 97.020 91.050 97.250 91.340 ;
        RECT 97.405 90.880 97.545 94.805 ;
        RECT 97.685 93.795 97.945 94.115 ;
        RECT 97.360 90.590 97.590 90.880 ;
        RECT 97.345 89.655 97.605 89.975 ;
        RECT 97.745 89.515 97.885 93.795 ;
        RECT 97.685 89.195 97.945 89.515 ;
        RECT 97.345 87.355 97.605 87.675 ;
        RECT 96.340 85.070 96.570 85.360 ;
        RECT 96.385 84.455 96.525 85.070 ;
        RECT 96.325 84.135 96.585 84.455 ;
        RECT 97.405 84.440 97.545 87.355 ;
        RECT 97.360 84.150 97.590 84.440 ;
        RECT 97.360 83.230 97.590 83.520 ;
        RECT 97.405 82.615 97.545 83.230 ;
        RECT 97.700 82.770 97.930 83.060 ;
        RECT 97.345 82.525 97.605 82.615 ;
        RECT 97.065 82.385 97.605 82.525 ;
        RECT 96.325 81.835 96.585 82.155 ;
        RECT 97.065 78.845 97.205 82.385 ;
        RECT 97.345 82.295 97.605 82.385 ;
        RECT 97.360 81.390 97.590 81.680 ;
        RECT 97.405 80.775 97.545 81.390 ;
        RECT 97.345 80.455 97.605 80.775 ;
        RECT 97.405 79.395 97.545 80.455 ;
        RECT 97.345 79.075 97.605 79.395 ;
        RECT 97.360 78.845 97.590 78.920 ;
        RECT 97.065 78.705 97.590 78.845 ;
        RECT 96.325 78.155 96.585 78.475 ;
        RECT 96.385 78.000 96.525 78.155 ;
        RECT 96.340 77.710 96.570 78.000 ;
        RECT 97.065 76.590 97.205 78.705 ;
        RECT 97.360 78.630 97.590 78.705 ;
        RECT 97.345 78.385 97.605 78.475 ;
        RECT 97.745 78.385 97.885 82.770 ;
        RECT 97.345 78.245 97.885 78.385 ;
        RECT 97.345 78.155 97.605 78.245 ;
        RECT 97.405 78.000 97.545 78.155 ;
        RECT 97.360 77.710 97.590 78.000 ;
        RECT 97.405 77.080 97.545 77.710 ;
        RECT 97.360 76.790 97.590 77.080 ;
        RECT 97.065 76.450 97.545 76.590 ;
        RECT 97.405 76.160 97.545 76.450 ;
        RECT 97.360 75.870 97.590 76.160 ;
        RECT 96.325 75.395 96.585 75.715 ;
        RECT 98.425 65.665 98.905 117.645 ;
        RECT 99.740 114.050 99.970 114.340 ;
        RECT 99.785 113.895 99.925 114.050 ;
        RECT 99.725 113.575 99.985 113.895 ;
        RECT 100.420 113.565 100.650 113.855 ;
        RECT 100.080 113.170 100.310 113.460 ;
        RECT 99.400 112.715 99.630 113.005 ;
        RECT 99.445 111.595 99.585 112.715 ;
        RECT 100.125 112.270 100.265 113.170 ;
        RECT 100.080 111.980 100.310 112.270 ;
        RECT 99.385 111.275 99.645 111.595 ;
        RECT 100.125 109.750 100.265 111.980 ;
        RECT 100.465 111.755 100.605 113.565 ;
        RECT 100.420 111.465 100.650 111.755 ;
        RECT 100.465 110.185 100.605 111.465 ;
        RECT 100.420 109.895 100.650 110.185 ;
        RECT 100.080 109.460 100.310 109.750 ;
        RECT 99.060 107.150 99.290 107.440 ;
        RECT 99.105 105.155 99.245 107.150 ;
        RECT 99.045 104.835 99.305 105.155 ;
        RECT 99.105 99.175 99.245 104.835 ;
        RECT 100.745 104.375 101.005 104.695 ;
        RECT 100.065 103.915 100.325 104.235 ;
        RECT 99.725 103.455 99.985 103.775 ;
        RECT 100.125 103.300 100.265 103.915 ;
        RECT 100.805 103.760 100.945 104.375 ;
        RECT 100.760 103.470 100.990 103.760 ;
        RECT 100.080 103.010 100.310 103.300 ;
        RECT 99.725 102.535 99.985 102.855 ;
        RECT 99.785 102.380 99.925 102.535 ;
        RECT 99.740 102.090 99.970 102.380 ;
        RECT 100.760 101.170 100.990 101.460 ;
        RECT 100.420 99.790 100.650 100.080 ;
        RECT 100.465 99.635 100.605 99.790 ;
        RECT 99.725 99.545 99.985 99.635 ;
        RECT 99.725 99.405 100.265 99.545 ;
        RECT 99.725 99.315 99.985 99.405 ;
        RECT 99.045 98.855 99.305 99.175 ;
        RECT 99.725 98.855 99.985 99.175 ;
        RECT 99.045 95.635 99.305 95.955 ;
        RECT 99.045 95.175 99.305 95.495 ;
        RECT 99.105 95.020 99.245 95.175 ;
        RECT 99.060 94.730 99.290 95.020 ;
        RECT 100.125 94.945 100.265 99.405 ;
        RECT 100.405 99.315 100.665 99.635 ;
        RECT 100.805 99.175 100.945 101.170 ;
        RECT 100.745 98.855 101.005 99.175 ;
        RECT 100.760 94.945 100.990 95.020 ;
        RECT 100.125 94.805 100.990 94.945 ;
        RECT 100.760 94.730 100.990 94.805 ;
        RECT 99.385 94.255 99.645 94.575 ;
        RECT 99.445 94.100 99.585 94.255 ;
        RECT 99.400 93.810 99.630 94.100 ;
        RECT 100.065 89.655 100.325 89.975 ;
        RECT 99.045 83.215 99.305 83.535 ;
        RECT 99.105 79.765 99.245 83.215 ;
        RECT 99.400 80.685 99.630 80.760 ;
        RECT 99.400 80.545 99.925 80.685 ;
        RECT 99.400 80.470 99.630 80.545 ;
        RECT 99.400 79.765 99.630 79.840 ;
        RECT 99.105 79.625 99.630 79.765 ;
        RECT 99.400 79.550 99.630 79.625 ;
        RECT 99.385 79.075 99.645 79.395 ;
        RECT 99.445 76.545 99.585 79.075 ;
        RECT 99.785 78.460 99.925 80.545 ;
        RECT 99.740 78.170 99.970 78.460 ;
        RECT 99.740 77.465 99.970 77.540 ;
        RECT 100.125 77.465 100.265 89.655 ;
        RECT 100.745 81.375 101.005 81.695 ;
        RECT 100.760 80.470 100.990 80.760 ;
        RECT 99.740 77.325 100.265 77.465 ;
        RECT 99.740 77.250 99.970 77.325 ;
        RECT 99.725 76.545 99.985 76.635 ;
        RECT 99.445 76.405 99.985 76.545 ;
        RECT 99.725 76.315 99.985 76.405 ;
        RECT 100.125 73.415 100.265 77.325 ;
        RECT 100.805 73.875 100.945 80.470 ;
        RECT 100.745 73.555 101.005 73.875 ;
        RECT 100.065 73.095 100.325 73.415 ;
        RECT 101.145 65.665 101.625 117.645 ;
        RECT 102.785 115.875 103.045 116.195 ;
        RECT 103.480 115.185 103.710 115.260 ;
        RECT 103.185 115.045 103.710 115.185 ;
        RECT 102.785 114.495 103.045 114.815 ;
        RECT 102.445 113.115 102.705 113.435 ;
        RECT 102.120 112.645 102.350 112.935 ;
        RECT 102.165 110.835 102.305 112.645 ;
        RECT 102.460 112.250 102.690 112.540 ;
        RECT 102.505 111.350 102.645 112.250 ;
        RECT 103.185 112.085 103.325 115.045 ;
        RECT 103.480 114.970 103.710 115.045 ;
        RECT 103.480 113.590 103.710 113.880 ;
        RECT 103.525 112.515 103.665 113.590 ;
        RECT 103.465 112.195 103.725 112.515 ;
        RECT 103.140 111.795 103.370 112.085 ;
        RECT 102.460 111.060 102.690 111.350 ;
        RECT 102.120 110.545 102.350 110.835 ;
        RECT 102.165 109.265 102.305 110.545 ;
        RECT 102.120 108.975 102.350 109.265 ;
        RECT 102.505 108.830 102.645 111.060 ;
        RECT 102.460 108.540 102.690 108.830 ;
        RECT 103.125 106.675 103.385 106.995 ;
        RECT 102.120 106.230 102.350 106.520 ;
        RECT 101.765 103.455 102.025 103.775 ;
        RECT 102.165 102.855 102.305 106.230 ;
        RECT 102.785 104.835 103.045 105.155 ;
        RECT 103.185 104.220 103.325 106.675 ;
        RECT 103.140 103.930 103.370 104.220 ;
        RECT 103.185 103.315 103.325 103.930 ;
        RECT 103.125 102.995 103.385 103.315 ;
        RECT 102.105 102.535 102.365 102.855 ;
        RECT 102.800 101.385 103.030 101.460 ;
        RECT 102.800 101.245 103.325 101.385 ;
        RECT 102.800 101.170 103.030 101.245 ;
        RECT 102.800 100.250 103.030 100.540 ;
        RECT 102.445 99.775 102.705 100.095 ;
        RECT 102.845 99.175 102.985 100.250 ;
        RECT 103.185 100.095 103.325 101.245 ;
        RECT 103.125 99.775 103.385 100.095 ;
        RECT 102.785 98.855 103.045 99.175 ;
        RECT 102.445 96.095 102.705 96.415 ;
        RECT 102.800 95.650 103.030 95.940 ;
        RECT 101.780 95.170 102.010 95.460 ;
        RECT 101.825 94.540 101.965 95.170 ;
        RECT 101.780 94.250 102.010 94.540 ;
        RECT 102.445 91.955 102.705 92.275 ;
        RECT 102.105 89.655 102.365 89.975 ;
        RECT 101.780 88.770 102.010 89.060 ;
        RECT 101.825 88.140 101.965 88.770 ;
        RECT 101.780 87.850 102.010 88.140 ;
        RECT 102.165 84.825 102.305 89.655 ;
        RECT 102.845 88.735 102.985 95.650 ;
        RECT 103.480 91.050 103.710 91.340 ;
        RECT 103.525 89.055 103.665 91.050 ;
        RECT 103.465 88.735 103.725 89.055 ;
        RECT 102.845 88.595 103.325 88.735 ;
        RECT 102.785 87.815 103.045 88.135 ;
        RECT 102.800 85.990 103.030 86.280 ;
        RECT 102.845 85.835 102.985 85.990 ;
        RECT 102.785 85.515 103.045 85.835 ;
        RECT 103.185 85.375 103.325 88.595 ;
        RECT 103.125 85.055 103.385 85.375 ;
        RECT 102.800 84.825 103.030 84.900 ;
        RECT 102.165 84.685 103.325 84.825 ;
        RECT 102.800 84.610 103.030 84.685 ;
        RECT 102.800 84.365 103.030 84.440 ;
        RECT 101.825 84.225 103.030 84.365 ;
        RECT 101.825 76.635 101.965 84.225 ;
        RECT 102.800 84.150 103.030 84.225 ;
        RECT 102.445 81.835 102.705 82.155 ;
        RECT 102.120 81.365 102.350 81.655 ;
        RECT 102.785 81.375 103.045 81.695 ;
        RECT 102.165 79.555 102.305 81.365 ;
        RECT 102.460 80.970 102.690 81.260 ;
        RECT 102.505 80.070 102.645 80.970 ;
        RECT 102.845 80.860 102.985 81.375 ;
        RECT 102.800 80.570 103.030 80.860 ;
        RECT 102.460 79.780 102.690 80.070 ;
        RECT 102.120 79.265 102.350 79.555 ;
        RECT 102.165 77.985 102.305 79.265 ;
        RECT 102.120 77.695 102.350 77.985 ;
        RECT 102.505 77.550 102.645 79.780 ;
        RECT 102.460 77.260 102.690 77.550 ;
        RECT 101.765 76.315 102.025 76.635 ;
        RECT 102.785 76.315 103.045 76.635 ;
        RECT 102.845 74.320 102.985 76.315 ;
        RECT 103.185 75.165 103.325 84.685 ;
        RECT 103.480 83.230 103.710 83.520 ;
        RECT 103.525 82.615 103.665 83.230 ;
        RECT 103.465 82.295 103.725 82.615 ;
        RECT 103.480 75.165 103.710 75.240 ;
        RECT 103.185 75.025 103.710 75.165 ;
        RECT 103.480 74.950 103.710 75.025 ;
        RECT 102.800 74.030 103.030 74.320 ;
        RECT 101.765 73.555 102.025 73.875 ;
        RECT 102.785 73.095 103.045 73.415 ;
        RECT 103.865 65.665 104.345 117.645 ;
        RECT 105.180 114.970 105.410 115.260 ;
        RECT 105.225 114.355 105.365 114.970 ;
        RECT 105.165 114.035 105.425 114.355 ;
        RECT 106.185 114.035 106.445 114.355 ;
        RECT 105.180 113.590 105.410 113.880 ;
        RECT 105.225 113.435 105.365 113.590 ;
        RECT 105.165 113.115 105.425 113.435 ;
        RECT 105.860 113.105 106.090 113.395 ;
        RECT 105.520 112.710 105.750 113.000 ;
        RECT 104.840 112.515 105.070 112.545 ;
        RECT 104.825 112.195 105.085 112.515 ;
        RECT 105.565 111.810 105.705 112.710 ;
        RECT 105.520 111.520 105.750 111.810 ;
        RECT 105.565 109.290 105.705 111.520 ;
        RECT 105.905 111.295 106.045 113.105 ;
        RECT 105.860 111.005 106.090 111.295 ;
        RECT 105.905 109.725 106.045 111.005 ;
        RECT 105.860 109.435 106.090 109.725 ;
        RECT 105.520 109.000 105.750 109.290 ;
        RECT 104.485 106.675 104.745 106.995 ;
        RECT 105.165 102.075 105.425 102.395 ;
        RECT 105.225 101.460 105.365 102.075 ;
        RECT 105.180 101.170 105.410 101.460 ;
        RECT 106.200 100.230 106.430 100.520 ;
        RECT 105.165 99.315 105.425 99.635 ;
        RECT 106.245 99.600 106.385 100.230 ;
        RECT 106.200 99.310 106.430 99.600 ;
        RECT 104.500 97.030 104.730 97.320 ;
        RECT 104.545 96.415 104.685 97.030 ;
        RECT 104.485 96.095 104.745 96.415 ;
        RECT 106.185 95.635 106.445 95.955 ;
        RECT 105.520 93.340 105.750 93.630 ;
        RECT 105.565 91.110 105.705 93.340 ;
        RECT 105.860 92.905 106.090 93.195 ;
        RECT 105.905 91.625 106.045 92.905 ;
        RECT 105.860 91.335 106.090 91.625 ;
        RECT 105.520 90.820 105.750 91.110 ;
        RECT 105.180 90.345 105.410 90.375 ;
        RECT 104.885 90.205 105.410 90.345 ;
        RECT 104.885 89.975 105.025 90.205 ;
        RECT 105.180 90.085 105.410 90.205 ;
        RECT 104.825 89.655 105.085 89.975 ;
        RECT 105.565 89.920 105.705 90.820 ;
        RECT 105.520 89.630 105.750 89.920 ;
        RECT 105.905 89.525 106.045 91.335 ;
        RECT 105.165 89.195 105.425 89.515 ;
        RECT 105.860 89.235 106.090 89.525 ;
        RECT 105.225 89.040 105.365 89.195 ;
        RECT 105.180 88.750 105.410 89.040 ;
        RECT 105.225 86.740 105.365 88.750 ;
        RECT 106.245 88.135 106.385 95.635 ;
        RECT 106.185 87.815 106.445 88.135 ;
        RECT 105.180 86.450 105.410 86.740 ;
        RECT 104.825 85.975 105.085 86.295 ;
        RECT 104.885 85.515 105.025 85.975 ;
        RECT 104.840 85.225 105.070 85.515 ;
        RECT 104.485 82.295 104.745 82.615 ;
        RECT 104.545 81.605 104.685 82.295 ;
        RECT 104.825 82.065 105.085 82.155 ;
        RECT 105.225 82.065 105.365 86.450 ;
        RECT 105.860 85.965 106.090 86.255 ;
        RECT 105.520 85.570 105.750 85.860 ;
        RECT 105.565 84.670 105.705 85.570 ;
        RECT 105.520 84.380 105.750 84.670 ;
        RECT 105.565 82.150 105.705 84.380 ;
        RECT 105.905 84.155 106.045 85.965 ;
        RECT 106.185 85.055 106.445 85.375 ;
        RECT 105.860 83.865 106.090 84.155 ;
        RECT 105.905 82.585 106.045 83.865 ;
        RECT 106.245 83.075 106.385 85.055 ;
        RECT 106.185 82.755 106.445 83.075 ;
        RECT 105.860 82.295 106.090 82.585 ;
        RECT 104.825 81.925 105.365 82.065 ;
        RECT 104.825 81.835 105.085 81.925 ;
        RECT 105.520 81.860 105.750 82.150 ;
        RECT 104.545 81.465 105.365 81.605 ;
        RECT 105.225 78.460 105.365 81.465 ;
        RECT 106.245 79.840 106.385 82.755 ;
        RECT 106.200 79.765 106.430 79.840 ;
        RECT 105.565 79.625 106.430 79.765 ;
        RECT 105.180 78.170 105.410 78.460 ;
        RECT 105.180 77.465 105.410 77.540 ;
        RECT 105.565 77.465 105.705 79.625 ;
        RECT 106.200 79.550 106.430 79.625 ;
        RECT 106.185 77.695 106.445 78.015 ;
        RECT 105.180 77.325 105.705 77.465 ;
        RECT 105.180 77.250 105.410 77.325 ;
        RECT 106.585 65.665 107.065 117.645 ;
        RECT 108.225 114.035 108.485 114.355 ;
        RECT 107.885 113.115 108.145 113.435 ;
        RECT 107.560 112.645 107.790 112.935 ;
        RECT 107.605 110.835 107.745 112.645 ;
        RECT 107.900 112.250 108.130 112.540 ;
        RECT 107.945 111.350 108.085 112.250 ;
        RECT 108.285 112.140 108.425 114.035 ;
        RECT 108.240 111.850 108.470 112.140 ;
        RECT 107.900 111.060 108.130 111.350 ;
        RECT 107.560 110.545 107.790 110.835 ;
        RECT 107.605 109.265 107.745 110.545 ;
        RECT 107.560 108.975 107.790 109.265 ;
        RECT 107.945 108.830 108.085 111.060 ;
        RECT 107.900 108.540 108.130 108.830 ;
        RECT 107.560 106.230 107.790 106.520 ;
        RECT 107.220 103.930 107.450 104.220 ;
        RECT 107.265 103.300 107.405 103.930 ;
        RECT 107.220 103.010 107.450 103.300 ;
        RECT 107.605 102.765 107.745 106.230 ;
        RECT 108.240 103.010 108.470 103.300 ;
        RECT 107.900 102.765 108.130 102.840 ;
        RECT 107.605 102.625 108.130 102.765 ;
        RECT 107.605 100.095 107.745 102.625 ;
        RECT 107.900 102.550 108.130 102.625 ;
        RECT 108.285 100.540 108.425 103.010 ;
        RECT 108.240 100.250 108.470 100.540 ;
        RECT 107.545 99.775 107.805 100.095 ;
        RECT 108.285 99.175 108.425 100.250 ;
        RECT 108.225 98.855 108.485 99.175 ;
        RECT 108.240 98.410 108.470 98.700 ;
        RECT 108.285 97.780 108.425 98.410 ;
        RECT 108.240 97.490 108.470 97.780 ;
        RECT 107.220 95.630 107.450 95.920 ;
        RECT 108.225 95.635 108.485 95.955 ;
        RECT 107.265 95.000 107.405 95.630 ;
        RECT 107.220 94.710 107.450 95.000 ;
        RECT 107.885 92.875 108.145 93.195 ;
        RECT 107.205 89.655 107.465 89.975 ;
        RECT 108.225 88.735 108.485 89.055 ;
        RECT 108.240 87.830 108.470 88.120 ;
        RECT 107.205 85.975 107.465 86.295 ;
        RECT 107.545 85.515 107.805 85.835 ;
        RECT 107.220 85.070 107.450 85.360 ;
        RECT 107.265 83.520 107.405 85.070 ;
        RECT 107.220 83.230 107.450 83.520 ;
        RECT 107.605 78.015 107.745 85.515 ;
        RECT 108.285 84.365 108.425 87.830 ;
        RECT 108.565 85.515 108.825 85.835 ;
        RECT 108.625 85.360 108.765 85.515 ;
        RECT 108.580 85.070 108.810 85.360 ;
        RECT 108.580 84.365 108.810 84.440 ;
        RECT 108.285 84.225 108.810 84.365 ;
        RECT 108.285 83.535 108.425 84.225 ;
        RECT 108.580 84.150 108.810 84.225 ;
        RECT 108.225 83.215 108.485 83.535 ;
        RECT 108.225 82.755 108.485 83.075 ;
        RECT 108.225 82.295 108.485 82.615 ;
        RECT 108.285 82.140 108.425 82.295 ;
        RECT 108.240 81.850 108.470 82.140 ;
        RECT 107.545 77.695 107.805 78.015 ;
        RECT 109.305 65.665 109.785 117.645 ;
        RECT 112.025 65.665 112.505 117.645 ;
        RECT 89.310 46.180 90.695 46.210 ;
        RECT 80.315 46.155 90.780 46.180 ;
        RECT 52.990 45.435 90.780 46.155 ;
        RECT 53.020 45.405 53.455 45.435 ;
        RECT 80.315 45.390 90.780 45.435 ;
        RECT 30.820 38.550 75.455 38.960 ;
        RECT 30.820 38.495 31.135 38.550 ;
        RECT 74.750 38.545 75.240 38.550 ;
        RECT 1.020 21.975 2.500 22.495 ;
        RECT 0.985 21.970 12.380 21.975 ;
        RECT 0.985 21.960 18.070 21.970 ;
        RECT 0.985 21.685 78.500 21.960 ;
        RECT 1.020 21.005 2.500 21.685 ;
        RECT 5.300 7.065 5.550 21.685 ;
        RECT 12.225 21.675 78.500 21.685 ;
        RECT 12.225 21.670 17.300 21.675 ;
        RECT 18.040 21.640 78.500 21.675 ;
        RECT 15.970 18.670 16.565 19.265 ;
        RECT 12.605 16.205 13.200 16.800 ;
        RECT 14.250 15.990 14.845 16.585 ;
        RECT 16.325 14.670 16.930 16.185 ;
        RECT 13.670 13.995 17.110 14.670 ;
        RECT 17.190 13.995 19.445 14.000 ;
        RECT 49.010 13.995 50.495 14.510 ;
        RECT 10.055 13.700 50.495 13.995 ;
        RECT 10.055 13.695 17.190 13.700 ;
        RECT 19.445 13.695 50.495 13.700 ;
        RECT 10.055 11.515 10.300 13.695 ;
        RECT 14.535 13.690 17.190 13.695 ;
        RECT 23.455 13.625 50.495 13.695 ;
        RECT 13.385 12.130 21.090 12.425 ;
        RECT 13.385 11.825 13.885 12.130 ;
        RECT 8.450 11.215 10.300 11.515 ;
        RECT 23.455 11.515 23.705 13.625 ;
        RECT 49.010 12.975 50.495 13.625 ;
        RECT 78.080 13.350 78.490 21.640 ;
        RECT 77.475 13.050 79.325 13.350 ;
        RECT 23.455 11.215 25.305 11.515 ;
        RECT 15.735 10.775 21.090 11.130 ;
        RECT 13.485 10.275 18.840 10.625 ;
        RECT 16.190 10.030 20.630 10.120 ;
        RECT 9.805 9.630 10.760 9.865 ;
        RECT 16.190 9.775 20.635 10.030 ;
        RECT 9.805 9.465 18.285 9.630 ;
        RECT 10.405 9.225 18.285 9.465 ;
        RECT 49.395 8.895 49.930 12.975 ;
        RECT 77.425 10.235 78.680 10.660 ;
        RECT 78.875 10.580 81.900 10.805 ;
        RECT 82.555 10.605 82.940 16.520 ;
        RECT 78.875 10.250 79.325 10.580 ;
        RECT 81.565 10.500 81.900 10.580 ;
        RECT 82.025 10.305 82.945 10.605 ;
        RECT 78.275 10.050 78.680 10.235 ;
        RECT 78.275 9.650 80.425 10.050 ;
        RECT 89.310 9.340 90.695 45.390 ;
        RECT 77.475 8.895 79.325 8.900 ;
        RECT 49.395 8.600 79.325 8.895 ;
        RECT 79.610 8.615 80.160 9.060 ;
        RECT 49.395 8.595 77.475 8.600 ;
        RECT 79.615 8.010 80.160 8.615 ;
        RECT 74.505 7.505 80.160 8.010 ;
        RECT 16.790 7.065 19.445 7.070 ;
        RECT 5.300 6.765 10.405 7.065 ;
        RECT 12.600 6.765 21.400 7.065 ;
        RECT 23.405 6.765 25.305 7.065 ;
        RECT 5.300 6.740 8.450 6.765 ;
        RECT 14.940 6.760 17.465 6.765 ;
        RECT 16.570 6.030 17.465 6.760 ;
        RECT 16.570 4.950 94.740 6.030 ;
        RECT 74.695 0.515 74.975 0.795 ;
        RECT 93.835 0.025 94.740 4.950 ;
      LAYER met2 ;
        RECT 55.505 225.200 55.785 225.480 ;
        RECT 58.275 225.200 58.555 225.480 ;
        RECT 61.015 225.185 61.295 225.465 ;
        RECT 63.785 225.200 64.065 225.480 ;
        RECT 66.525 225.210 66.805 225.490 ;
        RECT 69.330 225.235 69.610 225.515 ;
        RECT 48.990 204.000 50.490 204.205 ;
        RECT 48.990 203.315 50.495 204.000 ;
        RECT 48.990 203.195 50.490 203.315 ;
        RECT 78.275 116.105 78.595 116.165 ;
        RECT 80.995 116.105 81.315 116.165 ;
        RECT 78.275 115.965 81.315 116.105 ;
        RECT 78.275 115.905 78.595 115.965 ;
        RECT 80.995 115.905 81.315 115.965 ;
        RECT 97.315 116.105 97.635 116.165 ;
        RECT 102.755 116.105 103.075 116.165 ;
        RECT 97.315 115.965 103.075 116.105 ;
        RECT 97.315 115.905 97.635 115.965 ;
        RECT 102.755 115.905 103.075 115.965 ;
        RECT 78.955 115.645 79.275 115.705 ;
        RECT 88.815 115.645 89.135 115.705 ;
        RECT 91.875 115.645 92.195 115.705 ;
        RECT 107.660 115.645 108.030 115.715 ;
        RECT 78.955 115.505 89.135 115.645 ;
        RECT 78.955 115.445 79.275 115.505 ;
        RECT 88.815 115.445 89.135 115.505 ;
        RECT 89.415 115.505 108.030 115.645 ;
        RECT 69.775 115.185 70.095 115.245 ;
        RECT 72.495 115.185 72.815 115.245 ;
        RECT 80.460 115.185 80.830 115.255 ;
        RECT 89.415 115.185 89.555 115.505 ;
        RECT 91.875 115.445 92.195 115.505 ;
        RECT 107.660 115.435 108.030 115.505 ;
        RECT 69.775 115.045 80.830 115.185 ;
        RECT 69.775 114.985 70.095 115.045 ;
        RECT 72.495 114.985 72.815 115.045 ;
        RECT 80.460 114.975 80.830 115.045 ;
        RECT 84.135 115.045 89.555 115.185 ;
        RECT 69.095 114.725 69.415 114.785 ;
        RECT 73.660 114.725 74.030 114.795 ;
        RECT 69.095 114.585 74.030 114.725 ;
        RECT 69.095 114.525 69.415 114.585 ;
        RECT 73.660 114.515 74.030 114.585 ;
        RECT 61.615 114.265 61.935 114.325 ;
        RECT 74.535 114.265 74.855 114.325 ;
        RECT 61.615 114.125 74.855 114.265 ;
        RECT 61.615 114.065 61.935 114.125 ;
        RECT 74.535 114.065 74.855 114.125 ;
        RECT 77.595 114.265 77.915 114.325 ;
        RECT 84.135 114.265 84.275 115.045 ;
        RECT 89.155 114.725 89.475 114.785 ;
        RECT 91.875 114.725 92.195 114.785 ;
        RECT 89.155 114.585 92.195 114.725 ;
        RECT 89.155 114.525 89.475 114.585 ;
        RECT 91.875 114.525 92.195 114.585 ;
        RECT 96.295 114.725 96.615 114.785 ;
        RECT 100.860 114.725 101.230 114.795 ;
        RECT 102.755 114.725 103.075 114.785 ;
        RECT 96.295 114.585 103.075 114.725 ;
        RECT 96.295 114.525 96.615 114.585 ;
        RECT 100.860 114.515 101.230 114.585 ;
        RECT 102.755 114.525 103.075 114.585 ;
        RECT 77.595 114.125 84.275 114.265 ;
        RECT 94.060 114.265 94.430 114.335 ;
        RECT 96.975 114.265 97.295 114.325 ;
        RECT 105.135 114.265 105.455 114.325 ;
        RECT 94.060 114.125 105.455 114.265 ;
        RECT 77.595 114.065 77.915 114.125 ;
        RECT 94.060 114.055 94.430 114.125 ;
        RECT 96.975 114.065 97.295 114.125 ;
        RECT 105.135 114.065 105.455 114.125 ;
        RECT 106.155 114.265 106.475 114.325 ;
        RECT 108.195 114.265 108.515 114.325 ;
        RECT 106.155 114.125 108.515 114.265 ;
        RECT 106.155 114.065 106.475 114.125 ;
        RECT 108.195 114.065 108.515 114.125 ;
        RECT 66.860 113.865 67.230 113.875 ;
        RECT 66.860 113.805 67.375 113.865 ;
        RECT 70.115 113.805 70.435 113.865 ;
        RECT 66.860 113.665 70.435 113.805 ;
        RECT 66.860 113.605 67.375 113.665 ;
        RECT 70.115 113.605 70.435 113.665 ;
        RECT 77.060 113.805 77.430 113.875 ;
        RECT 77.935 113.805 78.255 113.865 ;
        RECT 80.995 113.805 81.315 113.865 ;
        RECT 77.060 113.665 81.315 113.805 ;
        RECT 66.860 113.595 67.230 113.605 ;
        RECT 77.060 113.595 77.430 113.665 ;
        RECT 77.935 113.605 78.255 113.665 ;
        RECT 80.995 113.605 81.315 113.665 ;
        RECT 83.860 113.805 84.230 113.875 ;
        RECT 97.315 113.805 97.635 113.865 ;
        RECT 99.695 113.805 100.015 113.865 ;
        RECT 83.860 113.665 97.635 113.805 ;
        RECT 83.860 113.595 84.230 113.665 ;
        RECT 97.315 113.605 97.635 113.665 ;
        RECT 99.615 113.605 100.015 113.805 ;
        RECT 61.955 113.345 62.275 113.405 ;
        RECT 64.675 113.345 64.995 113.405 ;
        RECT 61.955 113.205 64.995 113.345 ;
        RECT 61.955 113.145 62.275 113.205 ;
        RECT 64.675 113.145 64.995 113.205 ;
        RECT 70.115 113.345 70.435 113.405 ;
        RECT 75.895 113.345 76.215 113.405 ;
        RECT 83.375 113.345 83.695 113.405 ;
        RECT 70.115 113.205 76.215 113.345 ;
        RECT 70.115 113.145 70.435 113.205 ;
        RECT 75.895 113.145 76.215 113.205 ;
        RECT 81.085 113.205 83.695 113.345 ;
        RECT 81.085 112.945 81.225 113.205 ;
        RECT 83.375 113.145 83.695 113.205 ;
        RECT 92.555 113.345 92.875 113.405 ;
        RECT 94.935 113.345 95.255 113.405 ;
        RECT 99.615 113.345 99.755 113.605 ;
        RECT 102.415 113.345 102.735 113.405 ;
        RECT 105.135 113.345 105.455 113.405 ;
        RECT 107.855 113.345 108.175 113.405 ;
        RECT 92.555 113.205 108.175 113.345 ;
        RECT 92.555 113.145 92.875 113.205 ;
        RECT 94.935 113.145 95.255 113.205 ;
        RECT 102.415 113.145 102.735 113.205 ;
        RECT 105.135 113.145 105.455 113.205 ;
        RECT 107.855 113.145 108.175 113.205 ;
        RECT 65.015 112.885 65.335 112.945 ;
        RECT 66.375 112.885 66.695 112.945 ;
        RECT 65.015 112.745 66.695 112.885 ;
        RECT 65.015 112.685 65.335 112.745 ;
        RECT 66.375 112.685 66.695 112.745 ;
        RECT 72.495 112.885 72.815 112.945 ;
        RECT 75.215 112.885 75.535 112.945 ;
        RECT 72.495 112.745 75.535 112.885 ;
        RECT 72.495 112.685 72.815 112.745 ;
        RECT 75.215 112.685 75.535 112.745 ;
        RECT 80.995 112.685 81.315 112.945 ;
        RECT 65.355 112.425 65.675 112.485 ;
        RECT 67.055 112.425 67.375 112.485 ;
        RECT 72.495 112.425 72.815 112.485 ;
        RECT 81.085 112.425 81.225 112.685 ;
        RECT 65.355 112.285 81.225 112.425 ;
        RECT 81.675 112.425 81.995 112.485 ;
        RECT 83.035 112.425 83.355 112.485 ;
        RECT 81.675 112.285 83.355 112.425 ;
        RECT 65.355 112.225 65.675 112.285 ;
        RECT 67.055 112.225 67.375 112.285 ;
        RECT 72.495 112.225 72.815 112.285 ;
        RECT 81.675 112.225 81.995 112.285 ;
        RECT 83.035 112.225 83.355 112.285 ;
        RECT 103.435 112.425 103.755 112.485 ;
        RECT 104.795 112.425 105.115 112.485 ;
        RECT 103.435 112.285 105.115 112.425 ;
        RECT 103.435 112.225 103.755 112.285 ;
        RECT 104.795 112.225 105.115 112.285 ;
        RECT 70.795 111.965 71.115 112.025 ;
        RECT 75.555 111.965 75.875 112.025 ;
        RECT 70.795 111.825 75.875 111.965 ;
        RECT 70.795 111.765 71.115 111.825 ;
        RECT 75.555 111.765 75.875 111.825 ;
        RECT 74.535 111.505 74.855 111.565 ;
        RECT 77.255 111.505 77.575 111.565 ;
        RECT 74.535 111.365 77.575 111.505 ;
        RECT 74.535 111.305 74.855 111.365 ;
        RECT 77.255 111.305 77.575 111.365 ;
        RECT 97.995 111.505 98.315 111.565 ;
        RECT 99.355 111.505 99.675 111.565 ;
        RECT 97.995 111.365 99.675 111.505 ;
        RECT 97.995 111.305 98.315 111.365 ;
        RECT 99.355 111.305 99.675 111.365 ;
        RECT 67.055 111.045 67.375 111.105 ;
        RECT 69.095 111.045 69.415 111.105 ;
        RECT 67.055 110.905 69.415 111.045 ;
        RECT 67.055 110.845 67.375 110.905 ;
        RECT 69.095 110.845 69.415 110.905 ;
        RECT 75.555 111.045 75.875 111.105 ;
        RECT 96.295 111.045 96.615 111.105 ;
        RECT 75.555 110.905 96.615 111.045 ;
        RECT 75.555 110.845 75.875 110.905 ;
        RECT 96.295 110.845 96.615 110.905 ;
        RECT 70.260 109.205 70.630 109.275 ;
        RECT 77.935 109.205 78.255 109.265 ;
        RECT 70.260 109.065 78.255 109.205 ;
        RECT 70.260 108.995 70.630 109.065 ;
        RECT 77.935 109.005 78.255 109.065 ;
        RECT 88.815 109.205 89.135 109.265 ;
        RECT 104.260 109.205 104.630 109.275 ;
        RECT 88.815 109.065 104.630 109.205 ;
        RECT 88.815 109.005 89.135 109.065 ;
        RECT 104.260 108.995 104.630 109.065 ;
        RECT 75.895 108.745 76.215 108.805 ;
        RECT 90.660 108.745 91.030 108.815 ;
        RECT 97.315 108.745 97.635 108.805 ;
        RECT 75.895 108.605 84.275 108.745 ;
        RECT 75.895 108.545 76.215 108.605 ;
        RECT 84.135 108.285 84.275 108.605 ;
        RECT 90.660 108.605 97.635 108.745 ;
        RECT 90.660 108.535 91.030 108.605 ;
        RECT 97.315 108.545 97.635 108.605 ;
        RECT 97.460 108.285 97.830 108.355 ;
        RECT 84.135 108.145 97.830 108.285 ;
        RECT 97.460 108.075 97.830 108.145 ;
        RECT 103.095 106.905 103.415 106.965 ;
        RECT 104.455 106.905 104.775 106.965 ;
        RECT 103.095 106.765 104.775 106.905 ;
        RECT 103.095 106.705 103.415 106.765 ;
        RECT 104.455 106.705 104.775 106.765 ;
        RECT 62.635 106.445 62.955 106.505 ;
        RECT 68.075 106.445 68.395 106.505 ;
        RECT 70.115 106.445 70.435 106.505 ;
        RECT 62.635 106.305 70.435 106.445 ;
        RECT 62.635 106.245 62.955 106.305 ;
        RECT 68.075 106.245 68.395 106.305 ;
        RECT 70.115 106.245 70.435 106.305 ;
        RECT 84.395 106.445 84.715 106.505 ;
        RECT 86.775 106.445 87.095 106.505 ;
        RECT 91.875 106.445 92.195 106.505 ;
        RECT 84.395 106.305 92.195 106.445 ;
        RECT 84.395 106.245 84.715 106.305 ;
        RECT 86.775 106.245 87.095 106.305 ;
        RECT 91.875 106.245 92.195 106.305 ;
        RECT 86.095 105.985 86.415 106.045 ;
        RECT 88.475 105.985 88.795 106.045 ;
        RECT 90.855 105.985 91.175 106.045 ;
        RECT 86.095 105.845 91.175 105.985 ;
        RECT 86.095 105.785 86.415 105.845 ;
        RECT 88.475 105.785 88.795 105.845 ;
        RECT 90.855 105.785 91.175 105.845 ;
        RECT 86.435 105.065 86.755 105.125 ;
        RECT 88.135 105.065 88.455 105.125 ;
        RECT 88.815 105.065 89.135 105.125 ;
        RECT 84.655 104.925 89.135 105.065 ;
        RECT 63.995 103.685 64.315 103.745 ;
        RECT 67.395 103.685 67.715 103.745 ;
        RECT 70.115 103.685 70.435 103.745 ;
        RECT 63.995 103.545 70.435 103.685 ;
        RECT 63.995 103.485 64.315 103.545 ;
        RECT 67.395 103.485 67.715 103.545 ;
        RECT 70.115 103.485 70.435 103.545 ;
        RECT 80.995 103.685 81.315 103.745 ;
        RECT 83.715 103.685 84.035 103.745 ;
        RECT 84.655 103.685 84.795 104.925 ;
        RECT 86.435 104.865 86.755 104.925 ;
        RECT 88.135 104.865 88.455 104.925 ;
        RECT 88.815 104.865 89.135 104.925 ;
        RECT 99.015 105.065 99.335 105.125 ;
        RECT 102.755 105.065 103.075 105.125 ;
        RECT 99.015 104.925 103.075 105.065 ;
        RECT 99.015 104.865 99.335 104.925 ;
        RECT 102.755 104.865 103.075 104.925 ;
        RECT 96.975 104.605 97.295 104.665 ;
        RECT 100.715 104.605 101.035 104.665 ;
        RECT 96.975 104.465 101.035 104.605 ;
        RECT 96.975 104.405 97.295 104.465 ;
        RECT 100.715 104.405 101.035 104.465 ;
        RECT 87.115 104.145 87.435 104.205 ;
        RECT 91.535 104.145 91.855 104.205 ;
        RECT 94.255 104.145 94.575 104.205 ;
        RECT 97.315 104.145 97.635 104.205 ;
        RECT 100.035 104.145 100.355 104.205 ;
        RECT 87.115 104.005 100.355 104.145 ;
        RECT 87.115 103.945 87.435 104.005 ;
        RECT 91.535 103.945 91.855 104.005 ;
        RECT 94.255 103.945 94.575 104.005 ;
        RECT 97.315 103.945 97.635 104.005 ;
        RECT 100.035 103.945 100.355 104.005 ;
        RECT 85.415 103.685 85.735 103.745 ;
        RECT 80.995 103.545 84.795 103.685 ;
        RECT 80.995 103.485 81.315 103.545 ;
        RECT 83.715 103.485 84.035 103.545 ;
        RECT 85.335 103.485 85.735 103.685 ;
        RECT 88.135 103.685 88.455 103.745 ;
        RECT 90.855 103.685 91.175 103.745 ;
        RECT 95.275 103.685 95.595 103.745 ;
        RECT 96.975 103.685 97.295 103.745 ;
        RECT 88.135 103.545 97.295 103.685 ;
        RECT 88.135 103.485 88.455 103.545 ;
        RECT 90.855 103.485 91.175 103.545 ;
        RECT 95.275 103.485 95.595 103.545 ;
        RECT 96.975 103.485 97.295 103.545 ;
        RECT 99.695 103.685 100.015 103.745 ;
        RECT 101.735 103.685 102.055 103.745 ;
        RECT 99.695 103.545 102.055 103.685 ;
        RECT 99.695 103.485 100.015 103.545 ;
        RECT 101.735 103.485 102.055 103.545 ;
        RECT 62.635 102.765 62.955 102.825 ;
        RECT 66.715 102.765 67.035 102.825 ;
        RECT 70.115 102.765 70.435 102.825 ;
        RECT 71.815 102.765 72.135 102.825 ;
        RECT 62.635 102.625 64.395 102.765 ;
        RECT 62.635 102.565 62.955 102.625 ;
        RECT 64.255 102.365 64.395 102.625 ;
        RECT 66.715 102.625 72.135 102.765 ;
        RECT 66.715 102.565 67.035 102.625 ;
        RECT 70.115 102.565 70.435 102.625 ;
        RECT 71.815 102.565 72.135 102.625 ;
        RECT 79.975 102.765 80.295 102.825 ;
        RECT 83.375 102.765 83.695 102.825 ;
        RECT 85.335 102.765 85.475 103.485 ;
        RECT 97.655 103.225 97.975 103.285 ;
        RECT 103.095 103.225 103.415 103.285 ;
        RECT 97.575 103.085 103.415 103.225 ;
        RECT 97.575 103.025 97.975 103.085 ;
        RECT 103.095 103.025 103.415 103.085 ;
        RECT 88.815 102.765 89.135 102.825 ;
        RECT 89.835 102.765 90.155 102.825 ;
        RECT 79.975 102.625 90.155 102.765 ;
        RECT 79.975 102.565 80.295 102.625 ;
        RECT 83.375 102.565 83.695 102.625 ;
        RECT 88.815 102.565 89.135 102.625 ;
        RECT 89.835 102.565 90.155 102.625 ;
        RECT 94.595 102.765 94.915 102.825 ;
        RECT 97.575 102.765 97.715 103.025 ;
        RECT 94.595 102.625 97.715 102.765 ;
        RECT 99.695 102.765 100.015 102.825 ;
        RECT 102.075 102.765 102.395 102.825 ;
        RECT 99.695 102.625 102.475 102.765 ;
        RECT 94.595 102.565 94.915 102.625 ;
        RECT 99.695 102.565 100.015 102.625 ;
        RECT 102.075 102.565 102.475 102.625 ;
        RECT 63.120 100.385 63.490 102.265 ;
        RECT 64.255 102.165 64.655 102.365 ;
        RECT 64.335 102.105 64.655 102.165 ;
        RECT 65.015 102.305 65.335 102.365 ;
        RECT 66.715 102.305 67.035 102.365 ;
        RECT 65.015 102.165 67.035 102.305 ;
        RECT 102.335 102.305 102.475 102.565 ;
        RECT 105.135 102.305 105.455 102.365 ;
        RECT 65.015 102.105 65.335 102.165 ;
        RECT 66.715 102.105 67.035 102.165 ;
        RECT 68.560 100.385 68.930 102.265 ;
        RECT 70.115 100.465 70.435 100.525 ;
        RECT 69.695 100.325 73.745 100.465 ;
        RECT 74.000 100.385 74.370 102.265 ;
        RECT 79.440 100.385 79.810 102.265 ;
        RECT 84.880 100.385 85.250 102.265 ;
        RECT 88.135 101.385 88.455 101.445 ;
        RECT 88.815 101.385 89.135 101.445 ;
        RECT 88.135 101.245 89.135 101.385 ;
        RECT 88.135 101.185 88.455 101.245 ;
        RECT 88.815 101.185 89.135 101.245 ;
        RECT 90.320 100.385 90.690 102.265 ;
        RECT 95.760 100.385 96.130 102.265 ;
        RECT 101.200 100.385 101.570 102.265 ;
        RECT 102.335 102.165 105.455 102.305 ;
        RECT 105.135 102.105 105.455 102.165 ;
        RECT 106.640 100.385 107.010 102.265 ;
        RECT 112.080 100.385 112.450 102.265 ;
        RECT 61.615 100.005 61.935 100.065 ;
        RECT 65.015 100.005 65.335 100.065 ;
        RECT 61.615 99.865 65.335 100.005 ;
        RECT 61.615 99.805 61.935 99.865 ;
        RECT 65.015 99.805 65.335 99.865 ;
        RECT 68.075 100.005 68.395 100.065 ;
        RECT 69.695 100.005 69.835 100.325 ;
        RECT 70.115 100.265 70.435 100.325 ;
        RECT 68.075 99.865 69.835 100.005 ;
        RECT 70.115 100.005 70.435 100.065 ;
        RECT 72.495 100.005 72.815 100.065 ;
        RECT 70.115 99.865 72.815 100.005 ;
        RECT 73.605 100.005 73.745 100.325 ;
        RECT 80.995 100.005 81.315 100.065 ;
        RECT 83.375 100.005 83.695 100.065 ;
        RECT 73.605 99.865 83.695 100.005 ;
        RECT 68.075 99.805 68.395 99.865 ;
        RECT 70.115 99.805 70.435 99.865 ;
        RECT 72.495 99.805 72.815 99.865 ;
        RECT 80.995 99.805 81.315 99.865 ;
        RECT 83.295 99.805 83.695 99.865 ;
        RECT 84.055 100.005 84.375 100.065 ;
        RECT 86.095 100.005 86.415 100.065 ;
        RECT 84.055 99.865 86.415 100.005 ;
        RECT 84.055 99.805 84.375 99.865 ;
        RECT 86.095 99.805 86.415 99.865 ;
        RECT 86.775 100.005 87.095 100.065 ;
        RECT 102.415 100.005 102.735 100.065 ;
        RECT 86.775 99.865 102.735 100.005 ;
        RECT 86.775 99.805 87.095 99.865 ;
        RECT 102.415 99.805 102.735 99.865 ;
        RECT 103.095 100.005 103.415 100.065 ;
        RECT 107.515 100.005 107.835 100.065 ;
        RECT 103.095 99.865 107.835 100.005 ;
        RECT 103.095 99.805 103.415 99.865 ;
        RECT 107.515 99.805 107.835 99.865 ;
        RECT 83.295 99.545 83.435 99.805 ;
        RECT 88.135 99.545 88.455 99.605 ;
        RECT 83.295 99.405 88.455 99.545 ;
        RECT 88.135 99.345 88.455 99.405 ;
        RECT 90.855 99.545 91.175 99.605 ;
        RECT 93.575 99.545 93.895 99.605 ;
        RECT 90.855 99.405 93.895 99.545 ;
        RECT 90.855 99.345 91.175 99.405 ;
        RECT 93.575 99.345 93.895 99.405 ;
        RECT 94.255 99.545 94.575 99.605 ;
        RECT 95.275 99.545 95.595 99.605 ;
        RECT 97.315 99.545 97.635 99.605 ;
        RECT 99.695 99.545 100.015 99.605 ;
        RECT 94.255 99.405 100.015 99.545 ;
        RECT 94.255 99.345 94.575 99.405 ;
        RECT 95.275 99.345 95.595 99.405 ;
        RECT 97.315 99.345 97.635 99.405 ;
        RECT 99.695 99.345 100.015 99.405 ;
        RECT 100.375 99.545 100.695 99.605 ;
        RECT 105.135 99.545 105.455 99.605 ;
        RECT 100.375 99.405 105.455 99.545 ;
        RECT 100.375 99.345 100.695 99.405 ;
        RECT 105.135 99.345 105.455 99.405 ;
        RECT 69.095 99.085 69.415 99.145 ;
        RECT 75.895 99.085 76.215 99.145 ;
        RECT 69.095 98.945 76.215 99.085 ;
        RECT 69.095 98.885 69.415 98.945 ;
        RECT 67.395 98.625 67.715 98.685 ;
        RECT 69.435 98.625 69.755 98.685 ;
        RECT 60.400 96.685 60.770 98.565 ;
        RECT 61.615 97.245 61.935 97.305 ;
        RECT 63.655 97.245 63.975 97.305 ;
        RECT 61.615 97.105 63.975 97.245 ;
        RECT 61.615 97.045 61.935 97.105 ;
        RECT 63.655 97.045 63.975 97.105 ;
        RECT 65.840 96.685 66.210 98.565 ;
        RECT 67.395 98.485 69.755 98.625 ;
        RECT 67.395 98.425 67.715 98.485 ;
        RECT 69.435 98.425 69.755 98.485 ;
        RECT 69.775 98.165 70.095 98.225 ;
        RECT 70.545 98.165 70.685 98.945 ;
        RECT 75.895 98.885 76.215 98.945 ;
        RECT 81.675 99.085 81.995 99.145 ;
        RECT 86.435 99.085 86.755 99.145 ;
        RECT 81.675 98.945 86.755 99.085 ;
        RECT 81.675 98.885 81.995 98.945 ;
        RECT 86.435 98.885 86.755 98.945 ;
        RECT 87.115 99.085 87.435 99.145 ;
        RECT 91.875 99.085 92.195 99.145 ;
        RECT 87.115 98.945 92.195 99.085 ;
        RECT 87.115 98.885 87.435 98.945 ;
        RECT 91.875 98.885 92.195 98.945 ;
        RECT 96.975 99.085 97.295 99.145 ;
        RECT 99.015 99.085 99.335 99.145 ;
        RECT 99.695 99.085 100.015 99.145 ;
        RECT 96.975 98.945 100.015 99.085 ;
        RECT 96.975 98.885 97.295 98.945 ;
        RECT 99.015 98.885 99.335 98.945 ;
        RECT 99.695 98.885 100.015 98.945 ;
        RECT 100.715 99.085 101.035 99.145 ;
        RECT 102.755 99.085 103.075 99.145 ;
        RECT 108.195 99.085 108.515 99.145 ;
        RECT 100.715 98.945 108.515 99.085 ;
        RECT 100.715 98.885 101.035 98.945 ;
        RECT 102.755 98.885 103.075 98.945 ;
        RECT 108.195 98.885 108.515 98.945 ;
        RECT 88.135 98.625 88.455 98.685 ;
        RECT 88.815 98.625 89.135 98.685 ;
        RECT 69.775 98.025 70.685 98.165 ;
        RECT 69.775 97.965 70.095 98.025 ;
        RECT 71.280 96.685 71.650 98.565 ;
        RECT 76.720 96.685 77.090 98.565 ;
        RECT 82.160 96.685 82.530 98.565 ;
        RECT 83.375 96.785 83.695 96.845 ;
        RECT 83.295 96.585 83.695 96.785 ;
        RECT 84.395 96.785 84.715 96.845 ;
        RECT 86.435 96.785 86.755 96.845 ;
        RECT 84.395 96.645 86.755 96.785 ;
        RECT 87.600 96.685 87.970 98.565 ;
        RECT 88.135 98.485 89.135 98.625 ;
        RECT 88.135 98.425 88.455 98.485 ;
        RECT 88.815 98.425 89.135 98.485 ;
        RECT 88.815 98.165 89.135 98.225 ;
        RECT 92.555 98.165 92.875 98.225 ;
        RECT 88.815 98.025 92.875 98.165 ;
        RECT 88.815 97.965 89.135 98.025 ;
        RECT 90.775 97.765 90.915 98.025 ;
        RECT 92.555 97.965 92.875 98.025 ;
        RECT 90.775 97.565 91.175 97.765 ;
        RECT 90.855 97.505 91.175 97.565 ;
        RECT 88.815 97.045 89.135 97.305 ;
        RECT 88.905 96.785 89.045 97.045 ;
        RECT 91.875 96.785 92.195 96.845 ;
        RECT 88.905 96.645 92.195 96.785 ;
        RECT 93.040 96.685 93.410 98.565 ;
        RECT 98.480 96.685 98.850 98.565 ;
        RECT 103.920 96.685 104.290 98.565 ;
        RECT 109.360 96.685 109.730 98.565 ;
        RECT 84.395 96.585 84.715 96.645 ;
        RECT 86.435 96.585 86.755 96.645 ;
        RECT 91.875 96.585 92.195 96.645 ;
        RECT 62.635 96.325 62.955 96.385 ;
        RECT 66.375 96.325 66.695 96.385 ;
        RECT 62.635 96.185 66.695 96.325 ;
        RECT 62.635 96.125 62.955 96.185 ;
        RECT 66.375 96.125 66.695 96.185 ;
        RECT 70.795 96.325 71.115 96.385 ;
        RECT 83.295 96.325 83.435 96.585 ;
        RECT 70.795 96.185 83.435 96.325 ;
        RECT 102.415 96.325 102.735 96.385 ;
        RECT 104.455 96.325 104.775 96.385 ;
        RECT 102.415 96.185 104.775 96.325 ;
        RECT 70.795 96.125 71.115 96.185 ;
        RECT 102.415 96.125 102.735 96.185 ;
        RECT 104.455 96.125 104.775 96.185 ;
        RECT 64.335 95.865 64.655 95.925 ;
        RECT 69.095 95.865 69.415 95.925 ;
        RECT 64.335 95.725 69.415 95.865 ;
        RECT 64.335 95.665 64.655 95.725 ;
        RECT 69.095 95.665 69.415 95.725 ;
        RECT 70.115 95.865 70.435 95.925 ;
        RECT 72.835 95.865 73.155 95.925 ;
        RECT 83.375 95.865 83.695 95.925 ;
        RECT 70.115 95.665 70.515 95.865 ;
        RECT 72.835 95.725 83.695 95.865 ;
        RECT 72.835 95.665 73.155 95.725 ;
        RECT 83.375 95.665 83.695 95.725 ;
        RECT 91.535 95.865 91.855 95.925 ;
        RECT 99.015 95.865 99.335 95.925 ;
        RECT 91.535 95.725 99.335 95.865 ;
        RECT 91.535 95.665 91.855 95.725 ;
        RECT 99.015 95.665 99.335 95.725 ;
        RECT 106.155 95.865 106.475 95.925 ;
        RECT 108.195 95.865 108.515 95.925 ;
        RECT 106.155 95.725 108.515 95.865 ;
        RECT 106.155 95.665 106.475 95.725 ;
        RECT 108.195 95.665 108.515 95.725 ;
        RECT 67.395 95.405 67.715 95.465 ;
        RECT 69.775 95.405 70.095 95.465 ;
        RECT 67.395 95.265 70.095 95.405 ;
        RECT 70.375 95.405 70.515 95.665 ;
        RECT 70.795 95.405 71.115 95.465 ;
        RECT 70.375 95.265 71.115 95.405 ;
        RECT 67.395 95.205 67.715 95.265 ;
        RECT 69.775 95.205 70.095 95.265 ;
        RECT 70.795 95.205 71.115 95.265 ;
        RECT 81.675 95.405 81.995 95.465 ;
        RECT 85.415 95.405 85.735 95.465 ;
        RECT 81.675 95.265 85.735 95.405 ;
        RECT 81.675 95.205 81.995 95.265 ;
        RECT 85.415 95.205 85.735 95.265 ;
        RECT 94.595 95.405 94.915 95.465 ;
        RECT 96.635 95.405 96.955 95.465 ;
        RECT 99.015 95.405 99.335 95.465 ;
        RECT 94.595 95.265 99.335 95.405 ;
        RECT 94.595 95.205 94.915 95.265 ;
        RECT 96.635 95.205 96.955 95.265 ;
        RECT 99.015 95.205 99.335 95.265 ;
        RECT 86.435 94.945 86.755 95.005 ;
        RECT 96.975 94.945 97.295 95.005 ;
        RECT 83.295 94.805 86.755 94.945 ;
        RECT 64.335 94.485 64.655 94.545 ;
        RECT 66.375 94.485 66.695 94.545 ;
        RECT 64.335 94.345 66.695 94.485 ;
        RECT 64.335 94.285 64.655 94.345 ;
        RECT 66.375 94.285 66.695 94.345 ;
        RECT 68.075 94.485 68.395 94.545 ;
        RECT 83.295 94.485 83.435 94.805 ;
        RECT 86.435 94.745 86.755 94.805 ;
        RECT 92.815 94.805 97.295 94.945 ;
        RECT 68.075 94.345 83.435 94.485 ;
        RECT 83.860 94.485 84.230 94.555 ;
        RECT 92.815 94.485 92.955 94.805 ;
        RECT 96.975 94.745 97.295 94.805 ;
        RECT 83.860 94.345 92.955 94.485 ;
        RECT 93.575 94.485 93.895 94.545 ;
        RECT 99.355 94.485 99.675 94.545 ;
        RECT 93.575 94.345 99.675 94.485 ;
        RECT 68.075 94.285 68.395 94.345 ;
        RECT 83.860 94.275 84.230 94.345 ;
        RECT 93.575 94.285 93.895 94.345 ;
        RECT 99.355 94.285 99.675 94.345 ;
        RECT 63.995 94.025 64.315 94.085 ;
        RECT 66.375 94.025 66.695 94.085 ;
        RECT 63.995 93.885 66.695 94.025 ;
        RECT 63.995 93.825 64.315 93.885 ;
        RECT 66.375 93.825 66.695 93.885 ;
        RECT 81.675 94.025 81.995 94.085 ;
        RECT 88.135 94.025 88.455 94.085 ;
        RECT 81.675 93.885 88.455 94.025 ;
        RECT 81.675 93.825 81.995 93.885 ;
        RECT 88.135 93.825 88.455 93.885 ;
        RECT 89.835 94.025 90.155 94.085 ;
        RECT 90.855 94.025 91.175 94.085 ;
        RECT 89.835 93.885 91.175 94.025 ;
        RECT 89.835 93.825 90.155 93.885 ;
        RECT 90.855 93.825 91.175 93.885 ;
        RECT 95.275 94.025 95.595 94.085 ;
        RECT 97.655 94.025 97.975 94.085 ;
        RECT 95.275 93.885 97.975 94.025 ;
        RECT 95.275 93.825 95.595 93.885 ;
        RECT 97.655 93.825 97.975 93.885 ;
        RECT 61.955 93.565 62.275 93.625 ;
        RECT 68.075 93.565 68.395 93.625 ;
        RECT 61.955 93.425 68.395 93.565 ;
        RECT 61.955 93.365 62.275 93.425 ;
        RECT 68.075 93.365 68.395 93.425 ;
        RECT 81.335 93.565 81.655 93.625 ;
        RECT 86.775 93.565 87.095 93.625 ;
        RECT 89.155 93.565 89.475 93.625 ;
        RECT 81.335 93.425 89.475 93.565 ;
        RECT 81.335 93.365 81.655 93.425 ;
        RECT 86.775 93.365 87.095 93.425 ;
        RECT 89.155 93.365 89.475 93.425 ;
        RECT 90.855 93.565 91.175 93.625 ;
        RECT 96.975 93.565 97.295 93.625 ;
        RECT 90.855 93.425 97.295 93.565 ;
        RECT 90.855 93.365 91.175 93.425 ;
        RECT 96.975 93.365 97.295 93.425 ;
        RECT 79.975 93.105 80.295 93.165 ;
        RECT 89.835 93.105 90.155 93.165 ;
        RECT 79.975 92.965 90.155 93.105 ;
        RECT 79.975 92.905 80.295 92.965 ;
        RECT 89.835 92.905 90.155 92.965 ;
        RECT 91.535 93.105 91.855 93.165 ;
        RECT 107.855 93.105 108.175 93.165 ;
        RECT 91.535 92.965 108.175 93.105 ;
        RECT 91.535 92.905 91.855 92.965 ;
        RECT 107.855 92.905 108.175 92.965 ;
        RECT 66.715 92.645 67.035 92.705 ;
        RECT 72.835 92.645 73.155 92.705 ;
        RECT 77.935 92.645 78.255 92.705 ;
        RECT 66.715 92.505 78.255 92.645 ;
        RECT 66.715 92.445 67.035 92.505 ;
        RECT 72.835 92.445 73.155 92.505 ;
        RECT 77.935 92.445 78.255 92.505 ;
        RECT 80.655 92.645 80.975 92.705 ;
        RECT 83.375 92.645 83.695 92.705 ;
        RECT 80.655 92.505 83.695 92.645 ;
        RECT 80.655 92.445 80.975 92.505 ;
        RECT 83.375 92.445 83.695 92.505 ;
        RECT 88.815 92.645 89.135 92.705 ;
        RECT 90.855 92.645 91.175 92.705 ;
        RECT 88.815 92.505 91.175 92.645 ;
        RECT 88.815 92.445 89.135 92.505 ;
        RECT 90.855 92.445 91.175 92.505 ;
        RECT 83.860 92.245 84.230 92.255 ;
        RECT 76.235 92.185 76.555 92.245 ;
        RECT 83.035 92.185 83.355 92.245 ;
        RECT 76.235 92.045 83.355 92.185 ;
        RECT 76.235 91.985 76.555 92.045 ;
        RECT 83.035 91.985 83.355 92.045 ;
        RECT 83.715 91.985 84.230 92.245 ;
        RECT 89.835 92.185 90.155 92.245 ;
        RECT 102.415 92.185 102.735 92.245 ;
        RECT 89.835 92.045 102.735 92.185 ;
        RECT 89.835 91.985 90.155 92.045 ;
        RECT 102.415 91.985 102.735 92.045 ;
        RECT 83.860 91.975 84.230 91.985 ;
        RECT 81.675 91.725 81.995 91.785 ;
        RECT 86.580 91.725 86.950 91.795 ;
        RECT 46.840 91.585 86.950 91.725 ;
        RECT 46.840 91.580 81.995 91.585 ;
        RECT 46.840 22.515 47.480 91.580 ;
        RECT 81.675 91.525 81.995 91.580 ;
        RECT 86.580 91.515 86.950 91.585 ;
        RECT 64.140 91.265 64.510 91.335 ;
        RECT 86.435 91.265 86.755 91.325 ;
        RECT 47.990 91.125 86.755 91.265 ;
        RECT 47.990 91.115 64.510 91.125 ;
        RECT 0.995 21.005 2.485 22.505 ;
        RECT 46.790 20.785 47.495 22.515 ;
        RECT 11.310 20.260 47.460 20.785 ;
        RECT 11.310 16.800 11.805 20.260 ;
        RECT 47.995 19.940 48.480 91.115 ;
        RECT 64.140 91.055 64.510 91.115 ;
        RECT 86.435 91.065 86.755 91.125 ;
        RECT 65.015 90.805 65.335 90.865 ;
        RECT 67.055 90.805 67.375 90.865 ;
        RECT 62.215 90.665 67.375 90.805 ;
        RECT 61.615 90.345 61.935 90.405 ;
        RECT 62.215 90.345 62.355 90.665 ;
        RECT 65.015 90.605 65.335 90.665 ;
        RECT 67.055 90.605 67.375 90.665 ;
        RECT 77.935 90.805 78.255 90.865 ;
        RECT 81.675 90.805 81.995 90.865 ;
        RECT 77.935 90.665 81.995 90.805 ;
        RECT 77.935 90.605 78.255 90.665 ;
        RECT 81.675 90.605 81.995 90.665 ;
        RECT 61.615 90.205 62.355 90.345 ;
        RECT 87.115 90.345 87.435 90.405 ;
        RECT 88.815 90.345 89.135 90.405 ;
        RECT 87.115 90.205 89.135 90.345 ;
        RECT 61.615 90.145 61.935 90.205 ;
        RECT 87.115 90.145 87.435 90.205 ;
        RECT 88.815 90.145 89.135 90.205 ;
        RECT 70.795 89.885 71.115 89.945 ;
        RECT 74.535 89.885 74.855 89.945 ;
        RECT 70.795 89.745 74.855 89.885 ;
        RECT 70.795 89.685 71.115 89.745 ;
        RECT 74.535 89.685 74.855 89.745 ;
        RECT 82.695 89.885 83.015 89.945 ;
        RECT 97.315 89.885 97.635 89.945 ;
        RECT 100.035 89.885 100.355 89.945 ;
        RECT 102.075 89.885 102.395 89.945 ;
        RECT 82.695 89.745 102.395 89.885 ;
        RECT 82.695 89.685 83.015 89.745 ;
        RECT 97.315 89.685 97.635 89.745 ;
        RECT 100.035 89.685 100.355 89.745 ;
        RECT 102.075 89.685 102.395 89.745 ;
        RECT 104.795 89.885 105.115 89.945 ;
        RECT 107.175 89.885 107.495 89.945 ;
        RECT 104.795 89.745 107.495 89.885 ;
        RECT 104.795 89.685 105.115 89.745 ;
        RECT 107.175 89.685 107.495 89.745 ;
        RECT 97.655 89.425 97.975 89.485 ;
        RECT 105.135 89.425 105.455 89.485 ;
        RECT 97.655 89.285 105.455 89.425 ;
        RECT 97.655 89.225 97.975 89.285 ;
        RECT 105.135 89.225 105.455 89.285 ;
        RECT 67.735 88.965 68.055 89.025 ;
        RECT 75.895 88.965 76.215 89.025 ;
        RECT 67.735 88.825 76.215 88.965 ;
        RECT 67.735 88.765 68.055 88.825 ;
        RECT 75.895 88.765 76.215 88.825 ;
        RECT 103.435 88.965 103.755 89.025 ;
        RECT 108.195 88.965 108.515 89.025 ;
        RECT 103.435 88.825 108.515 88.965 ;
        RECT 103.435 88.765 103.755 88.825 ;
        RECT 108.195 88.765 108.515 88.825 ;
        RECT 72.495 88.505 72.815 88.565 ;
        RECT 87.115 88.505 87.435 88.565 ;
        RECT 93.915 88.505 94.235 88.565 ;
        RECT 72.495 88.365 94.235 88.505 ;
        RECT 72.495 88.305 72.815 88.365 ;
        RECT 87.115 88.305 87.435 88.365 ;
        RECT 93.915 88.305 94.235 88.365 ;
        RECT 65.355 88.045 65.675 88.105 ;
        RECT 70.455 88.045 70.775 88.105 ;
        RECT 71.815 88.045 72.135 88.105 ;
        RECT 65.355 87.905 72.135 88.045 ;
        RECT 65.355 87.845 65.675 87.905 ;
        RECT 70.455 87.845 70.775 87.905 ;
        RECT 71.815 87.845 72.135 87.905 ;
        RECT 83.715 88.045 84.035 88.105 ;
        RECT 88.815 88.045 89.135 88.105 ;
        RECT 83.715 87.905 89.135 88.045 ;
        RECT 83.715 87.845 84.035 87.905 ;
        RECT 88.815 87.845 89.135 87.905 ;
        RECT 102.755 88.045 103.075 88.105 ;
        RECT 106.155 88.045 106.475 88.105 ;
        RECT 102.755 87.905 106.475 88.045 ;
        RECT 102.755 87.845 103.075 87.905 ;
        RECT 106.155 87.845 106.475 87.905 ;
        RECT 66.375 87.585 66.695 87.645 ;
        RECT 67.055 87.585 67.375 87.645 ;
        RECT 66.375 87.445 67.375 87.585 ;
        RECT 66.375 87.385 66.695 87.445 ;
        RECT 67.055 87.385 67.375 87.445 ;
        RECT 91.195 87.585 91.515 87.645 ;
        RECT 93.575 87.585 93.895 87.645 ;
        RECT 97.315 87.585 97.635 87.645 ;
        RECT 91.195 87.445 97.635 87.585 ;
        RECT 91.195 87.385 91.515 87.445 ;
        RECT 93.575 87.385 93.895 87.445 ;
        RECT 97.315 87.385 97.635 87.445 ;
        RECT 68.075 87.125 68.395 87.185 ;
        RECT 73.515 87.125 73.835 87.185 ;
        RECT 68.075 86.985 73.835 87.125 ;
        RECT 68.075 86.925 68.395 86.985 ;
        RECT 73.515 86.925 73.835 86.985 ;
        RECT 78.275 86.665 78.595 86.725 ;
        RECT 80.995 86.665 81.315 86.725 ;
        RECT 78.275 86.525 81.315 86.665 ;
        RECT 78.275 86.465 78.595 86.525 ;
        RECT 80.995 86.465 81.315 86.525 ;
        RECT 70.115 86.205 70.435 86.265 ;
        RECT 71.815 86.205 72.135 86.265 ;
        RECT 70.115 86.065 72.135 86.205 ;
        RECT 70.115 86.005 70.435 86.065 ;
        RECT 71.815 86.005 72.135 86.065 ;
        RECT 104.795 86.205 105.115 86.265 ;
        RECT 107.175 86.205 107.495 86.265 ;
        RECT 104.795 86.065 107.495 86.205 ;
        RECT 104.795 86.005 105.115 86.065 ;
        RECT 107.175 86.005 107.495 86.065 ;
        RECT 102.755 85.745 103.075 85.805 ;
        RECT 107.515 85.745 107.835 85.805 ;
        RECT 108.535 85.745 108.855 85.805 ;
        RECT 102.755 85.605 108.855 85.745 ;
        RECT 102.755 85.545 103.075 85.605 ;
        RECT 107.515 85.545 107.835 85.605 ;
        RECT 108.535 85.545 108.855 85.605 ;
        RECT 68.075 85.285 68.395 85.345 ;
        RECT 71.815 85.285 72.135 85.345 ;
        RECT 68.075 85.145 72.135 85.285 ;
        RECT 68.075 85.085 68.395 85.145 ;
        RECT 71.815 85.085 72.135 85.145 ;
        RECT 89.495 85.285 89.815 85.345 ;
        RECT 92.215 85.285 92.535 85.345 ;
        RECT 89.495 85.145 92.535 85.285 ;
        RECT 89.495 85.085 89.815 85.145 ;
        RECT 92.215 85.085 92.535 85.145 ;
        RECT 103.095 85.285 103.415 85.345 ;
        RECT 106.155 85.285 106.475 85.345 ;
        RECT 103.095 85.145 106.475 85.285 ;
        RECT 103.095 85.085 103.415 85.145 ;
        RECT 106.155 85.085 106.475 85.145 ;
        RECT 92.555 84.365 92.875 84.425 ;
        RECT 96.295 84.365 96.615 84.425 ;
        RECT 92.555 84.225 96.615 84.365 ;
        RECT 92.555 84.165 92.875 84.225 ;
        RECT 96.295 84.165 96.615 84.225 ;
        RECT 72.155 83.905 72.475 83.965 ;
        RECT 77.595 83.905 77.915 83.965 ;
        RECT 72.155 83.765 77.915 83.905 ;
        RECT 72.155 83.705 72.475 83.765 ;
        RECT 77.595 83.705 77.915 83.765 ;
        RECT 66.715 83.445 67.035 83.505 ;
        RECT 69.435 83.445 69.755 83.505 ;
        RECT 72.495 83.445 72.815 83.505 ;
        RECT 66.715 83.305 72.815 83.445 ;
        RECT 66.715 83.245 67.035 83.305 ;
        RECT 69.435 83.245 69.755 83.305 ;
        RECT 72.495 83.245 72.815 83.305 ;
        RECT 92.555 83.445 92.875 83.505 ;
        RECT 93.915 83.445 94.235 83.505 ;
        RECT 99.015 83.445 99.335 83.505 ;
        RECT 108.195 83.445 108.515 83.505 ;
        RECT 92.555 83.305 94.235 83.445 ;
        RECT 92.555 83.245 92.875 83.305 ;
        RECT 93.915 83.245 94.235 83.305 ;
        RECT 94.855 83.305 108.515 83.445 ;
        RECT 65.355 82.985 65.675 83.045 ;
        RECT 67.055 82.985 67.375 83.045 ;
        RECT 72.155 82.985 72.475 83.045 ;
        RECT 65.355 82.845 72.475 82.985 ;
        RECT 65.355 82.785 65.675 82.845 ;
        RECT 67.055 82.785 67.375 82.845 ;
        RECT 72.155 82.785 72.475 82.845 ;
        RECT 92.215 82.985 92.535 83.045 ;
        RECT 94.855 82.985 94.995 83.305 ;
        RECT 99.015 83.245 99.335 83.305 ;
        RECT 108.195 83.245 108.515 83.305 ;
        RECT 92.215 82.845 94.995 82.985 ;
        RECT 106.155 82.985 106.475 83.045 ;
        RECT 108.195 82.985 108.515 83.045 ;
        RECT 106.155 82.845 108.515 82.985 ;
        RECT 92.215 82.785 92.535 82.845 ;
        RECT 106.155 82.785 106.475 82.845 ;
        RECT 108.195 82.785 108.515 82.845 ;
        RECT 66.375 82.525 66.695 82.585 ;
        RECT 71.815 82.525 72.135 82.585 ;
        RECT 64.255 82.385 72.135 82.525 ;
        RECT 61.955 82.065 62.275 82.125 ;
        RECT 63.655 82.065 63.975 82.125 ;
        RECT 64.255 82.065 64.395 82.385 ;
        RECT 66.375 82.325 66.695 82.385 ;
        RECT 71.815 82.325 72.135 82.385 ;
        RECT 92.215 82.525 92.535 82.585 ;
        RECT 95.275 82.525 95.595 82.585 ;
        RECT 97.315 82.525 97.635 82.585 ;
        RECT 92.215 82.385 97.635 82.525 ;
        RECT 92.215 82.325 92.535 82.385 ;
        RECT 95.275 82.325 95.595 82.385 ;
        RECT 97.315 82.325 97.635 82.385 ;
        RECT 103.435 82.525 103.755 82.585 ;
        RECT 104.455 82.525 104.775 82.585 ;
        RECT 108.195 82.525 108.515 82.585 ;
        RECT 103.435 82.385 108.515 82.525 ;
        RECT 103.435 82.325 103.755 82.385 ;
        RECT 104.455 82.325 104.775 82.385 ;
        RECT 108.195 82.325 108.515 82.385 ;
        RECT 61.955 81.925 64.395 82.065 ;
        RECT 70.115 82.065 70.435 82.125 ;
        RECT 80.655 82.065 80.975 82.125 ;
        RECT 70.115 81.925 80.975 82.065 ;
        RECT 61.955 81.865 62.275 81.925 ;
        RECT 63.655 81.865 63.975 81.925 ;
        RECT 70.115 81.865 70.435 81.925 ;
        RECT 80.655 81.865 80.975 81.925 ;
        RECT 90.855 82.065 91.175 82.125 ;
        RECT 96.295 82.065 96.615 82.125 ;
        RECT 102.415 82.065 102.735 82.125 ;
        RECT 104.795 82.065 105.115 82.125 ;
        RECT 90.855 81.925 96.615 82.065 ;
        RECT 90.855 81.865 91.175 81.925 ;
        RECT 96.295 81.865 96.615 81.925 ;
        RECT 97.745 81.925 105.115 82.065 ;
        RECT 67.055 81.605 67.375 81.665 ;
        RECT 70.795 81.605 71.115 81.665 ;
        RECT 72.155 81.605 72.475 81.665 ;
        RECT 67.055 81.465 72.475 81.605 ;
        RECT 67.055 81.405 67.375 81.465 ;
        RECT 70.795 81.405 71.115 81.465 ;
        RECT 72.155 81.405 72.475 81.465 ;
        RECT 87.115 81.605 87.435 81.665 ;
        RECT 89.155 81.605 89.475 81.665 ;
        RECT 92.215 81.605 92.535 81.665 ;
        RECT 87.115 81.465 92.535 81.605 ;
        RECT 87.115 81.405 87.435 81.465 ;
        RECT 89.155 81.405 89.475 81.465 ;
        RECT 92.215 81.405 92.535 81.465 ;
        RECT 70.795 81.145 71.115 81.205 ;
        RECT 71.815 81.145 72.135 81.205 ;
        RECT 70.795 81.005 72.135 81.145 ;
        RECT 70.795 80.945 71.115 81.005 ;
        RECT 71.815 80.945 72.135 81.005 ;
        RECT 78.615 81.145 78.935 81.205 ;
        RECT 81.335 81.145 81.655 81.205 ;
        RECT 83.375 81.145 83.695 81.205 ;
        RECT 85.755 81.145 86.075 81.205 ;
        RECT 78.615 81.005 86.075 81.145 ;
        RECT 78.615 80.945 78.935 81.005 ;
        RECT 81.335 80.945 81.655 81.005 ;
        RECT 83.375 80.945 83.695 81.005 ;
        RECT 85.755 80.945 86.075 81.005 ;
        RECT 94.255 81.145 94.575 81.205 ;
        RECT 97.745 81.145 97.885 81.925 ;
        RECT 102.415 81.865 102.735 81.925 ;
        RECT 104.795 81.865 105.115 81.925 ;
        RECT 100.715 81.605 101.035 81.665 ;
        RECT 102.755 81.605 103.075 81.665 ;
        RECT 100.715 81.465 103.075 81.605 ;
        RECT 100.715 81.405 101.035 81.465 ;
        RECT 102.755 81.405 103.075 81.465 ;
        RECT 94.255 81.005 97.885 81.145 ;
        RECT 94.255 80.945 94.575 81.005 ;
        RECT 75.895 80.685 76.215 80.745 ;
        RECT 77.255 80.685 77.575 80.745 ;
        RECT 75.895 80.545 77.575 80.685 ;
        RECT 75.895 80.485 76.215 80.545 ;
        RECT 77.255 80.485 77.575 80.545 ;
        RECT 79.975 80.685 80.295 80.745 ;
        RECT 83.375 80.685 83.695 80.745 ;
        RECT 86.095 80.685 86.415 80.745 ;
        RECT 79.975 80.545 86.415 80.685 ;
        RECT 79.975 80.485 80.295 80.545 ;
        RECT 83.375 80.485 83.695 80.545 ;
        RECT 86.095 80.485 86.415 80.545 ;
        RECT 92.555 80.685 92.875 80.745 ;
        RECT 97.315 80.685 97.635 80.745 ;
        RECT 92.555 80.545 97.635 80.685 ;
        RECT 92.555 80.485 92.875 80.545 ;
        RECT 97.315 80.485 97.635 80.545 ;
        RECT 62.635 80.225 62.955 80.285 ;
        RECT 64.675 80.225 64.995 80.285 ;
        RECT 62.635 80.085 64.995 80.225 ;
        RECT 62.635 80.025 62.955 80.085 ;
        RECT 64.675 80.025 64.995 80.085 ;
        RECT 68.075 80.225 68.395 80.285 ;
        RECT 72.495 80.225 72.815 80.285 ;
        RECT 75.215 80.225 75.535 80.285 ;
        RECT 81.335 80.225 81.655 80.285 ;
        RECT 82.695 80.225 83.015 80.285 ;
        RECT 87.115 80.225 87.435 80.285 ;
        RECT 68.075 80.085 87.435 80.225 ;
        RECT 68.075 80.025 68.395 80.085 ;
        RECT 72.495 80.025 72.815 80.085 ;
        RECT 75.215 80.025 75.535 80.085 ;
        RECT 81.335 80.025 81.655 80.085 ;
        RECT 82.695 80.025 83.015 80.085 ;
        RECT 87.115 80.025 87.435 80.085 ;
        RECT 75.895 79.765 76.215 79.825 ;
        RECT 78.615 79.765 78.935 79.825 ;
        RECT 87.115 79.765 87.435 79.825 ;
        RECT 88.475 79.765 88.795 79.825 ;
        RECT 75.895 79.625 78.935 79.765 ;
        RECT 75.895 79.565 76.215 79.625 ;
        RECT 78.615 79.565 78.935 79.625 ;
        RECT 84.135 79.625 88.795 79.765 ;
        RECT 77.255 79.305 77.575 79.365 ;
        RECT 84.135 79.305 84.275 79.625 ;
        RECT 87.115 79.565 87.435 79.625 ;
        RECT 88.475 79.565 88.795 79.625 ;
        RECT 77.255 79.165 84.275 79.305 ;
        RECT 97.315 79.305 97.635 79.365 ;
        RECT 99.355 79.305 99.675 79.365 ;
        RECT 97.315 79.165 99.675 79.305 ;
        RECT 77.255 79.105 77.575 79.165 ;
        RECT 97.315 79.105 97.635 79.165 ;
        RECT 99.355 79.105 99.675 79.165 ;
        RECT 78.955 78.845 79.275 78.905 ;
        RECT 79.975 78.845 80.295 78.905 ;
        RECT 78.955 78.705 80.295 78.845 ;
        RECT 78.955 78.645 79.275 78.705 ;
        RECT 79.975 78.645 80.295 78.705 ;
        RECT 89.155 78.845 89.475 78.905 ;
        RECT 89.155 78.705 97.545 78.845 ;
        RECT 89.155 78.645 89.475 78.705 ;
        RECT 97.405 78.445 97.545 78.705 ;
        RECT 78.275 78.385 78.595 78.445 ;
        RECT 80.315 78.385 80.635 78.445 ;
        RECT 83.375 78.385 83.695 78.445 ;
        RECT 78.275 78.245 83.695 78.385 ;
        RECT 78.275 78.185 78.595 78.245 ;
        RECT 80.315 78.185 80.635 78.245 ;
        RECT 83.375 78.185 83.695 78.245 ;
        RECT 90.855 78.385 91.175 78.445 ;
        RECT 96.295 78.385 96.615 78.445 ;
        RECT 90.855 78.245 96.615 78.385 ;
        RECT 90.855 78.185 91.175 78.245 ;
        RECT 96.295 78.185 96.615 78.245 ;
        RECT 97.315 78.185 97.635 78.445 ;
        RECT 84.395 77.925 84.715 77.985 ;
        RECT 86.775 77.925 87.095 77.985 ;
        RECT 84.395 77.785 87.095 77.925 ;
        RECT 84.395 77.725 84.715 77.785 ;
        RECT 86.775 77.725 87.095 77.785 ;
        RECT 89.155 77.925 89.475 77.985 ;
        RECT 94.255 77.925 94.575 77.985 ;
        RECT 89.155 77.785 94.575 77.925 ;
        RECT 89.155 77.725 89.475 77.785 ;
        RECT 94.255 77.725 94.575 77.785 ;
        RECT 106.155 77.925 106.475 77.985 ;
        RECT 107.515 77.925 107.835 77.985 ;
        RECT 106.155 77.785 107.835 77.925 ;
        RECT 106.155 77.725 106.475 77.785 ;
        RECT 107.515 77.725 107.835 77.785 ;
        RECT 92.555 77.465 92.875 77.525 ;
        RECT 93.915 77.465 94.235 77.525 ;
        RECT 92.555 77.325 94.235 77.465 ;
        RECT 92.555 77.265 92.875 77.325 ;
        RECT 93.915 77.265 94.235 77.325 ;
        RECT 78.955 77.005 79.275 77.065 ;
        RECT 80.995 77.005 81.315 77.065 ;
        RECT 78.955 76.865 81.315 77.005 ;
        RECT 78.955 76.805 79.275 76.865 ;
        RECT 80.995 76.805 81.315 76.865 ;
        RECT 83.375 76.545 83.695 76.605 ;
        RECT 85.415 76.545 85.735 76.605 ;
        RECT 83.375 76.405 85.735 76.545 ;
        RECT 83.375 76.345 83.695 76.405 ;
        RECT 85.415 76.345 85.735 76.405 ;
        RECT 86.775 76.545 87.095 76.605 ;
        RECT 88.135 76.545 88.455 76.605 ;
        RECT 86.775 76.405 88.455 76.545 ;
        RECT 86.775 76.345 87.095 76.405 ;
        RECT 88.135 76.345 88.455 76.405 ;
        RECT 99.695 76.545 100.015 76.605 ;
        RECT 101.735 76.545 102.055 76.605 ;
        RECT 102.755 76.545 103.075 76.605 ;
        RECT 99.695 76.405 103.075 76.545 ;
        RECT 99.695 76.345 100.015 76.405 ;
        RECT 101.735 76.345 102.055 76.405 ;
        RECT 102.755 76.345 103.075 76.405 ;
        RECT 69.095 76.085 69.415 76.145 ;
        RECT 70.115 76.085 70.435 76.145 ;
        RECT 69.095 75.945 70.435 76.085 ;
        RECT 69.095 75.885 69.415 75.945 ;
        RECT 70.115 75.885 70.435 75.945 ;
        RECT 92.215 75.625 92.535 75.685 ;
        RECT 96.295 75.625 96.615 75.685 ;
        RECT 92.215 75.485 96.615 75.625 ;
        RECT 92.215 75.425 92.535 75.485 ;
        RECT 96.295 75.425 96.615 75.485 ;
        RECT 62.295 75.165 62.615 75.225 ;
        RECT 70.455 75.165 70.775 75.225 ;
        RECT 77.255 75.165 77.575 75.225 ;
        RECT 62.295 75.025 77.575 75.165 ;
        RECT 62.295 74.965 62.615 75.025 ;
        RECT 70.455 74.965 70.775 75.025 ;
        RECT 77.255 74.965 77.575 75.025 ;
        RECT 86.775 74.705 87.095 74.765 ;
        RECT 88.135 74.705 88.455 74.765 ;
        RECT 86.775 74.565 88.455 74.705 ;
        RECT 86.775 74.505 87.095 74.565 ;
        RECT 88.135 74.505 88.455 74.565 ;
        RECT 81.675 73.785 81.995 73.845 ;
        RECT 86.435 73.785 86.755 73.845 ;
        RECT 81.675 73.645 86.755 73.785 ;
        RECT 81.675 73.585 81.995 73.645 ;
        RECT 86.435 73.585 86.755 73.645 ;
        RECT 100.715 73.785 101.035 73.845 ;
        RECT 101.735 73.785 102.055 73.845 ;
        RECT 100.715 73.645 102.055 73.785 ;
        RECT 100.715 73.585 101.035 73.645 ;
        RECT 101.735 73.585 102.055 73.645 ;
        RECT 69.095 73.325 69.415 73.385 ;
        RECT 71.815 73.325 72.135 73.385 ;
        RECT 69.095 73.185 72.135 73.325 ;
        RECT 69.095 73.125 69.415 73.185 ;
        RECT 71.815 73.125 72.135 73.185 ;
        RECT 100.035 73.325 100.355 73.385 ;
        RECT 102.755 73.325 103.075 73.385 ;
        RECT 100.035 73.185 103.075 73.325 ;
        RECT 100.035 73.125 100.355 73.185 ;
        RECT 102.755 73.125 103.075 73.185 ;
        RECT 63.120 70.385 63.490 72.265 ;
        RECT 68.560 70.385 68.930 72.265 ;
        RECT 74.000 70.385 74.370 72.265 ;
        RECT 79.440 70.385 79.810 72.265 ;
        RECT 84.880 70.385 85.250 72.265 ;
        RECT 90.320 70.385 90.690 72.265 ;
        RECT 95.760 70.385 96.130 72.265 ;
        RECT 101.200 70.385 101.570 72.265 ;
        RECT 106.640 70.385 107.010 72.265 ;
        RECT 112.080 70.385 112.450 72.265 ;
        RECT 60.400 66.685 60.770 68.565 ;
        RECT 65.840 66.685 66.210 68.565 ;
        RECT 71.280 66.685 71.650 68.565 ;
        RECT 76.720 66.685 77.090 68.565 ;
        RECT 82.160 66.685 82.530 68.565 ;
        RECT 87.600 66.685 87.970 68.565 ;
        RECT 93.040 66.685 93.410 68.565 ;
        RECT 98.480 66.685 98.850 68.565 ;
        RECT 103.920 66.685 104.290 68.565 ;
        RECT 109.360 66.685 109.730 68.565 ;
        RECT 74.750 38.545 75.240 38.955 ;
        RECT 15.970 19.255 75.425 19.265 ;
        RECT 15.970 18.645 152.700 19.255 ;
        RECT 74.540 18.635 152.700 18.645 ;
        RECT 75.425 18.560 152.700 18.635 ;
        RECT 11.310 16.205 13.200 16.800 ;
        RECT 14.250 16.475 56.115 16.505 ;
        RECT 56.120 16.475 133.385 16.515 ;
        RECT 11.310 15.495 11.805 16.205 ;
        RECT 14.250 15.990 133.385 16.475 ;
        RECT 55.210 15.985 133.385 15.990 ;
        RECT 55.545 15.980 133.385 15.985 ;
        RECT 56.120 15.975 133.385 15.980 ;
        RECT 6.985 14.975 11.805 15.495 ;
        RECT 6.985 4.520 7.505 14.975 ;
        RECT 11.310 14.970 11.805 14.975 ;
        RECT 49.000 12.995 50.490 14.495 ;
        RECT 15.730 10.780 48.455 11.130 ;
        RECT 15.730 10.775 16.135 10.780 ;
        RECT 77.430 10.245 90.690 10.670 ;
        RECT 74.655 7.590 74.935 7.870 ;
        RECT 9.710 6.765 24.115 7.070 ;
        RECT 6.985 4.515 112.980 4.520 ;
        RECT 6.985 4.005 114.090 4.515 ;
        RECT 6.985 3.995 35.650 4.005 ;
        RECT 36.770 3.995 114.090 4.005 ;
        RECT 7.515 3.990 35.650 3.995 ;
        RECT 74.695 0.515 74.975 0.795 ;
        RECT 94.100 0.405 94.380 0.685 ;
        RECT 113.180 0.000 114.085 3.995 ;
        RECT 132.495 -0.010 133.385 15.975 ;
        RECT 151.810 0.010 152.700 18.560 ;
      LAYER met3 ;
        RECT 54.980 224.235 56.480 225.745 ;
        RECT 57.750 224.235 59.250 225.745 ;
        RECT 60.490 224.220 61.990 225.730 ;
        RECT 63.260 224.235 64.760 225.745 ;
        RECT 66.000 224.245 67.500 225.755 ;
        RECT 68.805 224.270 70.305 225.780 ;
        RECT 103.315 206.170 118.315 207.170 ;
        RECT 100.315 205.170 110.315 206.170 ;
        RECT 111.315 205.170 122.315 206.170 ;
        RECT 48.990 204.005 50.490 204.200 ;
        RECT 97.315 204.170 102.315 205.170 ;
        RECT 119.315 204.170 124.315 205.170 ;
        RECT 48.990 203.310 50.495 204.005 ;
        RECT 48.990 203.190 50.490 203.310 ;
        RECT 95.315 203.170 99.315 204.170 ;
        RECT 122.315 203.170 126.315 204.170 ;
        RECT 93.315 202.170 97.315 203.170 ;
        RECT 124.315 202.170 128.315 203.170 ;
        RECT 91.315 201.170 95.315 202.170 ;
        RECT 126.315 201.170 130.315 202.170 ;
        RECT 90.315 200.170 93.315 201.170 ;
        RECT 128.315 200.170 131.315 201.170 ;
        RECT 89.315 199.170 92.315 200.170 ;
        RECT 130.315 199.170 133.315 200.170 ;
        RECT 88.315 198.170 90.315 199.170 ;
        RECT 131.315 198.170 134.315 199.170 ;
        RECT 87.315 197.170 89.315 198.170 ;
        RECT 132.315 197.170 135.315 198.170 ;
        RECT 86.315 196.170 88.315 197.170 ;
        RECT 133.315 196.170 136.315 197.170 ;
        RECT 85.315 195.170 87.315 196.170 ;
        RECT 134.315 195.170 137.315 196.170 ;
        RECT 84.315 194.170 86.315 195.170 ;
        RECT 135.315 194.170 137.315 195.170 ;
        RECT 83.315 193.170 85.315 194.170 ;
        RECT 136.315 193.170 138.315 194.170 ;
        RECT 82.315 192.170 85.315 193.170 ;
        RECT 82.315 191.170 84.315 192.170 ;
        RECT 99.315 191.170 123.315 193.170 ;
        RECT 137.315 192.170 139.315 193.170 ;
        RECT 137.315 191.170 140.315 192.170 ;
        RECT 81.315 190.170 83.315 191.170 ;
        RECT 80.315 189.170 83.315 190.170 ;
        RECT 100.315 189.170 122.315 191.170 ;
        RECT 138.315 190.170 140.315 191.170 ;
        RECT 80.315 188.170 82.315 189.170 ;
        RECT 101.315 188.170 121.315 189.170 ;
        RECT 139.315 188.170 141.315 190.170 ;
        RECT 79.315 185.170 81.315 188.170 ;
        RECT 101.315 187.170 120.315 188.170 ;
        RECT 102.315 186.170 120.315 187.170 ;
        RECT 140.315 186.170 142.315 188.170 ;
        RECT 78.315 183.170 80.315 185.170 ;
        RECT 103.315 184.170 119.315 186.170 ;
        RECT 78.315 182.170 79.315 183.170 ;
        RECT 96.315 182.170 97.315 183.170 ;
        RECT 104.315 182.170 118.315 184.170 ;
        RECT 141.315 183.170 143.315 186.170 ;
        RECT 125.315 182.170 126.315 183.170 ;
        RECT 77.315 178.170 79.315 182.170 ;
        RECT 95.315 180.170 98.315 182.170 ;
        RECT 105.315 181.170 117.315 182.170 ;
        RECT 105.315 180.170 116.315 181.170 ;
        RECT 124.315 180.170 127.315 182.170 ;
        RECT 142.315 180.170 144.315 183.170 ;
        RECT 94.315 178.170 99.315 180.170 ;
        RECT 106.315 179.170 116.315 180.170 ;
        RECT 77.315 175.170 78.315 178.170 ;
        RECT 93.315 177.170 100.315 178.170 ;
        RECT 107.315 177.170 115.315 179.170 ;
        RECT 123.315 178.170 128.315 180.170 ;
        RECT 143.315 179.170 144.315 180.170 ;
        RECT 122.315 177.170 129.315 178.170 ;
        RECT 92.315 175.170 101.315 177.170 ;
        RECT 108.315 175.170 114.315 177.170 ;
        RECT 121.315 176.170 129.315 177.170 ;
        RECT 121.315 175.170 130.315 176.170 ;
        RECT 76.315 172.170 78.315 175.170 ;
        RECT 91.315 173.170 102.315 175.170 ;
        RECT 109.315 174.170 113.315 175.170 ;
        RECT 90.315 172.170 103.315 173.170 ;
        RECT 110.315 172.170 112.315 174.170 ;
        RECT 120.315 173.170 131.315 175.170 ;
        RECT 77.315 169.170 78.315 172.170 ;
        RECT 89.315 171.170 103.315 172.170 ;
        RECT 119.315 171.170 132.315 173.170 ;
        RECT 89.315 170.170 104.315 171.170 ;
        RECT 118.315 170.170 133.315 171.170 ;
        RECT 77.315 165.170 79.315 169.170 ;
        RECT 88.315 168.170 105.315 170.170 ;
        RECT 117.315 168.170 134.315 170.170 ;
        RECT 143.315 168.170 145.315 179.170 ;
        RECT 87.315 166.170 106.315 168.170 ;
        RECT 116.315 166.170 135.315 168.170 ;
        RECT 143.315 167.170 144.315 168.170 ;
        RECT 86.315 165.170 107.315 166.170 ;
        RECT 115.315 165.170 136.315 166.170 ;
        RECT 78.315 164.170 79.315 165.170 ;
        RECT 85.315 164.170 107.315 165.170 ;
        RECT 114.315 164.170 136.315 165.170 ;
        RECT 142.315 164.170 144.315 167.170 ;
        RECT 78.315 162.170 80.315 164.170 ;
        RECT 85.315 163.170 108.315 164.170 ;
        RECT 114.315 163.170 137.315 164.170 ;
        RECT 79.315 159.170 81.315 162.170 ;
        RECT 84.315 161.170 109.315 163.170 ;
        RECT 113.315 161.170 138.315 163.170 ;
        RECT 141.315 161.170 143.315 164.170 ;
        RECT 140.315 159.170 142.315 161.170 ;
        RECT 80.315 157.170 82.315 159.170 ;
        RECT 139.315 157.170 141.315 159.170 ;
        RECT 81.315 156.170 83.315 157.170 ;
        RECT 82.315 154.170 84.315 156.170 ;
        RECT 138.315 155.170 140.315 157.170 ;
        RECT 137.315 154.170 139.315 155.170 ;
        RECT 83.315 153.170 85.315 154.170 ;
        RECT 136.315 153.170 138.315 154.170 ;
        RECT 84.315 152.170 86.315 153.170 ;
        RECT 135.315 152.170 137.315 153.170 ;
        RECT 85.315 151.170 87.315 152.170 ;
        RECT 134.315 151.170 137.315 152.170 ;
        RECT 85.315 150.170 88.315 151.170 ;
        RECT 133.315 150.170 136.315 151.170 ;
        RECT 86.315 149.170 89.315 150.170 ;
        RECT 132.315 149.170 135.315 150.170 ;
        RECT 88.315 148.170 90.315 149.170 ;
        RECT 131.315 148.170 134.315 149.170 ;
        RECT 89.315 147.170 92.315 148.170 ;
        RECT 130.315 147.170 133.315 148.170 ;
        RECT 90.315 146.170 93.315 147.170 ;
        RECT 128.315 146.170 131.315 147.170 ;
        RECT 91.315 145.170 95.315 146.170 ;
        RECT 127.315 145.170 130.315 146.170 ;
        RECT 93.315 144.170 97.315 145.170 ;
        RECT 124.315 144.170 128.315 145.170 ;
        RECT 95.315 143.170 99.315 144.170 ;
        RECT 122.315 143.170 127.315 144.170 ;
        RECT 97.315 142.170 102.315 143.170 ;
        RECT 119.315 142.170 124.315 143.170 ;
        RECT 99.315 141.170 108.315 142.170 ;
        RECT 114.315 141.170 122.315 142.170 ;
        RECT 103.315 140.170 118.315 141.170 ;
        RECT 67.345 120.280 70.145 122.785 ;
        RECT 70.745 120.280 73.545 122.785 ;
        RECT 74.145 120.280 76.945 122.785 ;
        RECT 77.545 120.280 80.345 122.785 ;
        RECT 80.945 120.280 83.745 122.785 ;
        RECT 91.145 119.730 93.945 122.970 ;
        RECT 94.545 119.730 97.345 122.970 ;
        RECT 97.945 119.730 100.745 122.970 ;
        RECT 101.345 119.730 104.145 122.970 ;
        RECT 104.745 119.730 107.545 122.970 ;
        RECT 63.495 107.215 63.795 119.165 ;
        RECT 66.895 113.900 67.195 119.165 ;
        RECT 66.880 113.570 67.210 113.900 ;
        RECT 70.295 109.300 70.595 119.165 ;
        RECT 73.695 114.820 73.995 119.165 ;
        RECT 73.680 114.490 74.010 114.820 ;
        RECT 77.095 113.900 77.395 119.165 ;
        RECT 80.495 115.280 80.795 119.165 ;
        RECT 80.480 114.950 80.810 115.280 ;
        RECT 83.895 113.900 84.195 119.165 ;
        RECT 77.080 113.570 77.410 113.900 ;
        RECT 83.880 113.570 84.210 113.900 ;
        RECT 70.280 108.970 70.610 109.300 ;
        RECT 87.295 107.215 87.595 119.165 ;
        RECT 90.695 108.840 90.995 119.165 ;
        RECT 94.095 114.360 94.395 119.165 ;
        RECT 94.080 114.030 94.410 114.360 ;
        RECT 90.680 108.510 91.010 108.840 ;
        RECT 97.495 108.380 97.795 119.165 ;
        RECT 100.895 114.820 101.195 119.165 ;
        RECT 100.880 114.490 101.210 114.820 ;
        RECT 104.295 109.300 104.595 119.165 ;
        RECT 107.695 115.740 107.995 119.165 ;
        RECT 107.680 115.410 108.010 115.740 ;
        RECT 104.280 108.970 104.610 109.300 ;
        RECT 97.480 108.050 97.810 108.380 ;
        RECT 63.495 106.915 64.475 107.215 ;
        RECT 1.010 100.300 60.005 102.325 ;
        RECT 63.140 100.335 63.470 102.315 ;
        RECT 52.045 72.350 53.990 100.300 ;
        RECT 60.420 96.635 60.750 98.615 ;
        RECT 64.175 91.360 64.475 106.915 ;
        RECT 86.615 106.915 87.595 107.215 ;
        RECT 68.580 100.335 68.910 102.315 ;
        RECT 74.020 100.335 74.350 102.315 ;
        RECT 79.460 100.335 79.790 102.315 ;
        RECT 84.900 100.335 85.230 102.315 ;
        RECT 65.860 96.635 66.190 98.615 ;
        RECT 71.300 96.635 71.630 98.615 ;
        RECT 76.740 96.635 77.070 98.615 ;
        RECT 82.180 96.635 82.510 98.615 ;
        RECT 83.880 94.250 84.210 94.580 ;
        RECT 83.895 92.280 84.195 94.250 ;
        RECT 83.880 91.950 84.210 92.280 ;
        RECT 86.615 91.820 86.915 106.915 ;
        RECT 90.340 100.335 90.670 102.315 ;
        RECT 95.780 100.335 96.110 102.315 ;
        RECT 101.220 100.335 101.550 102.315 ;
        RECT 106.660 100.335 106.990 102.315 ;
        RECT 112.100 100.335 112.430 102.315 ;
        RECT 87.620 96.635 87.950 98.615 ;
        RECT 93.060 96.635 93.390 98.615 ;
        RECT 98.500 96.635 98.830 98.615 ;
        RECT 103.940 96.635 104.270 98.615 ;
        RECT 109.380 96.635 109.710 98.615 ;
        RECT 86.600 91.490 86.930 91.820 ;
        RECT 64.160 91.030 64.490 91.360 ;
        RECT 52.005 70.325 61.830 72.350 ;
        RECT 63.140 70.335 63.470 72.315 ;
        RECT 68.580 70.335 68.910 72.315 ;
        RECT 74.020 70.335 74.350 72.315 ;
        RECT 79.460 70.335 79.790 72.315 ;
        RECT 84.900 70.335 85.230 72.315 ;
        RECT 90.340 70.335 90.670 72.315 ;
        RECT 95.780 70.335 96.110 72.315 ;
        RECT 101.220 70.335 101.550 72.315 ;
        RECT 106.660 70.335 106.990 72.315 ;
        RECT 112.100 70.335 112.430 72.315 ;
        RECT 52.045 70.305 53.990 70.325 ;
        RECT 60.420 66.635 60.750 68.615 ;
        RECT 65.860 66.635 66.190 68.615 ;
        RECT 71.300 66.635 71.630 68.615 ;
        RECT 76.740 66.635 77.070 68.615 ;
        RECT 82.180 66.635 82.510 68.615 ;
        RECT 87.620 66.635 87.950 68.615 ;
        RECT 93.060 66.635 93.390 68.615 ;
        RECT 98.500 66.635 98.830 68.615 ;
        RECT 103.940 66.635 104.270 68.615 ;
        RECT 109.380 66.635 109.710 68.615 ;
        RECT 1.000 20.995 2.500 22.505 ;
        RECT 47.995 10.780 48.460 20.990 ;
        RECT 49.005 12.985 50.505 14.495 ;
        RECT 74.495 1.625 75.450 38.975 ;
        RECT 74.170 0.160 75.670 1.625 ;
        RECT 74.170 0.020 75.685 0.160 ;
        RECT 93.575 0.005 95.075 1.515 ;
        RECT 112.945 0.000 114.445 1.510 ;
        RECT 132.265 -0.010 133.765 1.500 ;
        RECT 151.575 0.010 153.075 1.520 ;
      LAYER met4 ;
        RECT 66.510 225.765 66.865 225.780 ;
        RECT 58.260 225.755 58.595 225.760 ;
        RECT 54.985 224.230 56.485 225.745 ;
        RECT 57.745 224.230 59.255 225.755 ;
        RECT 60.485 224.220 61.990 225.760 ;
        RECT 63.240 224.230 64.755 225.740 ;
        RECT 66.010 224.240 67.480 225.765 ;
        RECT 68.800 224.270 70.310 225.780 ;
        RECT 48.995 133.650 49.000 135.660 ;
        RECT 50.500 133.650 51.005 135.660 ;
        RECT 50.500 120.235 70.320 122.735 ;
        RECT 79.795 120.270 94.345 122.770 ;
        RECT 55.935 100.325 60.345 102.325 ;
        RECT 55.935 100.320 60.840 100.325 ;
        RECT 50.500 98.625 62.345 98.640 ;
        RECT 50.500 96.625 60.345 98.625 ;
        RECT 50.500 96.575 62.345 96.625 ;
        RECT 55.975 72.325 60.380 72.350 ;
        RECT 55.975 70.325 112.505 72.325 ;
        RECT 50.500 66.640 112.505 68.625 ;
        RECT 60.345 66.625 112.505 66.640 ;
        RECT 50.500 55.235 50.525 56.730 ;
        RECT 48.995 31.160 49.000 32.655 ;
        RECT 74.160 -0.010 75.690 1.615 ;
        RECT 93.530 0.000 95.030 1.520 ;
        RECT 112.925 0.000 114.450 1.495 ;
        RECT 132.225 0.035 133.785 1.495 ;
        RECT 132.490 0.000 133.385 0.035 ;
        RECT 151.570 0.005 153.075 1.515 ;
      LAYER met5 ;
        RECT 76.235 100.615 78.235 102.035 ;
        RECT 106.235 100.615 108.235 102.035 ;
        RECT 79.935 96.915 81.935 98.335 ;
        RECT 109.935 96.915 111.935 98.335 ;
        RECT 76.235 70.615 78.235 72.035 ;
        RECT 106.235 70.615 108.235 72.035 ;
        RECT 79.935 66.915 81.935 68.335 ;
        RECT 109.935 66.915 111.935 68.335 ;
  END
END tt_um_vco_mix_dac
END LIBRARY

